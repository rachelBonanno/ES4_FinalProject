library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity background_rom is
  port(
	  clk : in std_logic;
	  row_idx: in unsigned(6 downto 0);
	  col_idx : in unsigned(5 downto 0); 
	  rgb : out std_logic_vector(5 downto 0)
	  );
end background_rom;

architecture synth of background_rom is

signal location : std_logic_vector(12 downto 0);
begin
	process (clk) begin
		if rising_edge(clk) then
			case location is
			
				when "0000010010100" => rgb <= "100001";
				when "0000010010101" => rgb <= "100001";
				when "0000010010110" => rgb <= "100001";
				when "0000010010111" => rgb <= "100001";
				when "0000010011000" => rgb <= "100001";
				when "0000010011001" => rgb <= "100001";
				when "0000010011010" => rgb <= "100001";
				when "0000010011101" => rgb <= "100001";
				when "0000010011110" => rgb <= "100001";
				when "0000010100010" => rgb <= "100001";
				when "0000010100011" => rgb <= "100001";
				when "0000010100110" => rgb <= "100001";
				when "0000010100111" => rgb <= "100001";
				when "0000010101000" => rgb <= "100001";
				when "0000010101001" => rgb <= "100001";
				when "0000010101101" => rgb <= "100001";
				when "0000010101110" => rgb <= "100001";
				when "0000010110000" => rgb <= "100001";
				when "0000010110001" => rgb <= "100001";
				when "0000010110010" => rgb <= "100001";
				when "0000010110110" => rgb <= "100001";
				when "0000010110111" => rgb <= "100001";
				when "0000010111000" => rgb <= "100001";
				when "0000010111001" => rgb <= "100001";
				when "0000100010100" => rgb <= "100001";
				when "0000100010101" => rgb <= "100001";
				when "0000100010110" => rgb <= "100001";
				when "0000100010111" => rgb <= "100001";
				when "0000100011000" => rgb <= "100001";
				when "0000100011001" => rgb <= "100001";
				when "0000100011010" => rgb <= "100001";
				when "0000100011101" => rgb <= "100001";
				when "0000100011110" => rgb <= "100001";
				when "0000100100010" => rgb <= "100001";
				when "0000100100011" => rgb <= "100001";
				when "0000100100110" => rgb <= "100001";
				when "0000100100111" => rgb <= "100001";
				when "0000100101000" => rgb <= "100001";
				when "0000100101001" => rgb <= "100001";
				when "0000100101101" => rgb <= "100001";
				when "0000100101110" => rgb <= "100001";
				when "0000100101111" => rgb <= "100001";
				when "0000100110000" => rgb <= "100001";
				when "0000100110001" => rgb <= "100001";
				when "0000100110110" => rgb <= "100001";
				when "0000100110111" => rgb <= "100001";
				when "0000100111000" => rgb <= "100001";
				when "0000100111001" => rgb <= "100001";
				when "0000110010111" => rgb <= "100001";
				when "0000110011000" => rgb <= "100001";
				when "0000110011101" => rgb <= "100001";
				when "0000110011110" => rgb <= "100001";
				when "0000110100010" => rgb <= "100001";
				when "0000110100011" => rgb <= "100001";
				when "0000110100110" => rgb <= "100001";
				when "0000110100111" => rgb <= "100001";
				when "0000110101101" => rgb <= "100001";
				when "0000110101110" => rgb <= "100001";
				when "0000110101111" => rgb <= "100001";
				when "0000110110000" => rgb <= "100001";
				when "0000110110110" => rgb <= "100001";
				when "0000110110111" => rgb <= "100001";
				when "0001000010111" => rgb <= "100001";
				when "0001000011000" => rgb <= "100001";
				when "0001000011101" => rgb <= "100001";
				when "0001000011110" => rgb <= "100001";
				when "0001000100010" => rgb <= "100001";
				when "0001000100011" => rgb <= "100001";
				when "0001000100110" => rgb <= "100001";
				when "0001000100111" => rgb <= "100001";
				when "0001000101000" => rgb <= "100001";
				when "0001000101001" => rgb <= "100001";
				when "0001000101101" => rgb <= "100001";
				when "0001000101110" => rgb <= "100001";
				when "0001000101111" => rgb <= "100001";
				when "0001000110000" => rgb <= "100001";
				when "0001000110110" => rgb <= "100001";
				when "0001000110111" => rgb <= "100001";
				when "0001000111000" => rgb <= "100001";
				when "0001000111001" => rgb <= "100001";
				when "0001010010111" => rgb <= "100001";
				when "0001010011000" => rgb <= "100001";
				when "0001010011101" => rgb <= "100001";
				when "0001010011110" => rgb <= "100001";
				when "0001010100010" => rgb <= "100001";
				when "0001010100011" => rgb <= "100001";
				when "0001010101000" => rgb <= "100001";
				when "0001010101001" => rgb <= "100001";
				when "0001010101101" => rgb <= "100001";
				when "0001010101110" => rgb <= "100001";
				when "0001010101111" => rgb <= "100001";
				when "0001010110000" => rgb <= "100001";
				when "0001010110001" => rgb <= "100001";
				when "0001010111000" => rgb <= "100001";
				when "0001010111001" => rgb <= "100001";
				when "0001100010111" => rgb <= "100001";
				when "0001100011000" => rgb <= "100001";
				when "0001100011101" => rgb <= "100001";
				when "0001100011110" => rgb <= "100001";
				when "0001100011111" => rgb <= "100001";
				when "0001100100000" => rgb <= "100001";
				when "0001100100001" => rgb <= "100001";
				when "0001100100010" => rgb <= "100001";
				when "0001100100011" => rgb <= "100001";
				when "0001100100110" => rgb <= "100001";
				when "0001100100111" => rgb <= "100001";
				when "0001100101000" => rgb <= "100001";
				when "0001100101001" => rgb <= "100001";
				when "0001100101101" => rgb <= "100001";
				when "0001100101110" => rgb <= "100001";
				when "0001100101111" => rgb <= "100001";
				when "0001100110000" => rgb <= "100001";
				when "0001100110001" => rgb <= "100001";
				when "0001100110010" => rgb <= "100001";
				when "0001100110110" => rgb <= "100001";
				when "0001100110111" => rgb <= "100001";
				when "0001100111000" => rgb <= "100001";
				when "0001100111001" => rgb <= "100001";
				when "0001110010111" => rgb <= "100001";
				when "0001110011000" => rgb <= "100001";
				when "0001110011110" => rgb <= "100001";
				when "0001110011111" => rgb <= "100001";
				when "0001110100000" => rgb <= "100001";
				when "0001110100001" => rgb <= "100001";
				when "0001110100010" => rgb <= "100001";
				when "0001110100110" => rgb <= "100001";
				when "0001110100111" => rgb <= "100001";
				when "0001110101000" => rgb <= "100001";
				when "0001110101001" => rgb <= "100001";
				when "0001110101101" => rgb <= "100001";
				when "0001110101110" => rgb <= "100001";
				when "0001110110000" => rgb <= "100001";
				when "0001110110001" => rgb <= "100001";
				when "0001110110010" => rgb <= "100001";
				when "0001110110110" => rgb <= "100001";
				when "0001110110111" => rgb <= "100001";
				when "0001110111000" => rgb <= "100001";
				when "0001110111001" => rgb <= "100001";
				when "0010100000001" => rgb <= "111111";
				when "0010100000010" => rgb <= "111111";
				when "0010100000011" => rgb <= "111111";
				when "0010100000101" => rgb <= "111111";
				when "0010100001000" => rgb <= "111111";
				when "0010100001001" => rgb <= "111111";
				when "0010100001010" => rgb <= "111111";
				when "0010100001100" => rgb <= "111111";
				when "0010100001110" => rgb <= "111111";
				when "0010100010000" => rgb <= "111111";
				when "0010100010001" => rgb <= "111111";
				when "0010100010011" => rgb <= "111111";
				when "0010100010100" => rgb <= "111111";
				when "0010100010101" => rgb <= "111111";
				when "0010100011000" => rgb <= "111111";
				when "0010100011001" => rgb <= "111111";
				when "0010100110101" => rgb <= "111111";
				when "0010100110110" => rgb <= "111111";
				when "0010100110111" => rgb <= "111111";
				when "0010100111001" => rgb <= "111111";
				when "0010100111100" => rgb <= "111111";
				when "0010100111101" => rgb <= "111111";
				when "0010100111110" => rgb <= "111111";
				when "0010101000000" => rgb <= "111111";
				when "0010101000010" => rgb <= "111111";
				when "0010101000100" => rgb <= "111111";
				when "0010101000101" => rgb <= "111111";
				when "0010101000111" => rgb <= "111111";
				when "0010101001000" => rgb <= "111111";
				when "0010101001001" => rgb <= "111111";
				when "0010101001100" => rgb <= "111111";
				when "0010101001101" => rgb <= "111111";
				when "0010110000001" => rgb <= "111111";
				when "0010110000011" => rgb <= "111111";
				when "0010110000101" => rgb <= "111111";
				when "0010110001000" => rgb <= "111111";
				when "0010110001010" => rgb <= "111111";
				when "0010110001100" => rgb <= "111111";
				when "0010110001110" => rgb <= "111111";
				when "0010110010000" => rgb <= "111111";
				when "0010110010011" => rgb <= "111111";
				when "0010110010101" => rgb <= "111111";
				when "0010110011001" => rgb <= "111111";
				when "0010110110101" => rgb <= "111111";
				when "0010110110111" => rgb <= "111111";
				when "0010110111001" => rgb <= "111111";
				when "0010110111100" => rgb <= "111111";
				when "0010110111110" => rgb <= "111111";
				when "0010111000000" => rgb <= "111111";
				when "0010111000010" => rgb <= "111111";
				when "0010111000100" => rgb <= "111111";
				when "0010111000111" => rgb <= "111111";
				when "0010111001001" => rgb <= "111111";
				when "0010111001011" => rgb <= "111111";
				when "0010111001110" => rgb <= "111111";
				when "0011000000001" => rgb <= "111111";
				when "0011000000010" => rgb <= "111111";
				when "0011000000011" => rgb <= "111111";
				when "0011000000101" => rgb <= "111111";
				when "0011000001000" => rgb <= "111111";
				when "0011000001001" => rgb <= "111111";
				when "0011000001010" => rgb <= "111111";
				when "0011000001101" => rgb <= "111111";
				when "0011000010000" => rgb <= "111111";
				when "0011000010001" => rgb <= "111111";
				when "0011000010011" => rgb <= "111111";
				when "0011000010100" => rgb <= "111111";
				when "0011000010101" => rgb <= "111111";
				when "0011000011001" => rgb <= "111111";
				when "0011000110101" => rgb <= "111111";
				when "0011000110110" => rgb <= "111111";
				when "0011000110111" => rgb <= "111111";
				when "0011000111001" => rgb <= "111111";
				when "0011000111100" => rgb <= "111111";
				when "0011000111101" => rgb <= "111111";
				when "0011000111110" => rgb <= "111111";
				when "0011001000001" => rgb <= "111111";
				when "0011001000100" => rgb <= "111111";
				when "0011001000101" => rgb <= "111111";
				when "0011001000111" => rgb <= "111111";
				when "0011001001000" => rgb <= "111111";
				when "0011001001001" => rgb <= "111111";
				when "0011001001101" => rgb <= "111111";
				when "0011001001110" => rgb <= "111111";
				when "0011010000001" => rgb <= "111111";
				when "0011010000101" => rgb <= "111111";
				when "0011010001000" => rgb <= "111111";
				when "0011010001010" => rgb <= "111111";
				when "0011010001101" => rgb <= "111111";
				when "0011010010000" => rgb <= "111111";
				when "0011010010011" => rgb <= "111111";
				when "0011010010100" => rgb <= "111111";
				when "0011010011001" => rgb <= "111111";
				when "0011010110101" => rgb <= "111111";
				when "0011010111001" => rgb <= "111111";
				when "0011010111100" => rgb <= "111111";
				when "0011010111110" => rgb <= "111111";
				when "0011011000001" => rgb <= "111111";
				when "0011011000100" => rgb <= "111111";
				when "0011011000111" => rgb <= "111111";
				when "0011011001000" => rgb <= "111111";
				when "0011011001100" => rgb <= "111111";
				when "0011100000001" => rgb <= "111111";
				when "0011100000101" => rgb <= "111111";
				when "0011100000110" => rgb <= "111111";
				when "0011100001000" => rgb <= "111111";
				when "0011100001010" => rgb <= "111111";
				when "0011100001101" => rgb <= "111111";
				when "0011100010000" => rgb <= "111111";
				when "0011100010001" => rgb <= "111111";
				when "0011100010011" => rgb <= "111111";
				when "0011100010101" => rgb <= "111111";
				when "0011100011000" => rgb <= "111111";
				when "0011100011001" => rgb <= "111111";
				when "0011100011010" => rgb <= "111111";
				when "0011100110101" => rgb <= "111111";
				when "0011100111001" => rgb <= "111111";
				when "0011100111010" => rgb <= "111111";
				when "0011100111100" => rgb <= "111111";
				when "0011100111110" => rgb <= "111111";
				when "0011101000001" => rgb <= "111111";
				when "0011101000100" => rgb <= "111111";
				when "0011101000101" => rgb <= "111111";
				when "0011101000111" => rgb <= "111111";
				when "0011101001001" => rgb <= "111111";
				when "0011101001100" => rgb <= "111111";
				when "0011101001101" => rgb <= "111111";
				when "0011101001110" => rgb <= "111111";
				when "1000000011000" => rgb <= "111111";
				when "1000000011001" => rgb <= "111111";
				when "1000000011010" => rgb <= "111111";
				when "1000000011011" => rgb <= "111111";
				when "1000000011100" => rgb <= "111111";
				when "1000000011101" => rgb <= "111111";
				when "1000000011110" => rgb <= "111111";
				when "1000000011111" => rgb <= "111111";
				when "1000000100000" => rgb <= "111111";
				when "1000000100001" => rgb <= "111111";
				when "1000000100010" => rgb <= "111111";
				when "1000000100011" => rgb <= "111111";
				when "1000000100100" => rgb <= "111111";
				when "1000000100101" => rgb <= "111111";
				when "1000000100110" => rgb <= "111111";
				when "1000000100111" => rgb <= "111111";
				when "1000000101000" => rgb <= "111111";
				when "1000000101001" => rgb <= "111111";
				when "1000000101010" => rgb <= "111111";
				when "1000000101011" => rgb <= "111111";
				when "1000000101100" => rgb <= "111111";
				when "1000000101101" => rgb <= "111111";
				when "1000000101110" => rgb <= "111111";
				when "1000000101111" => rgb <= "111111";
				when "1000000110000" => rgb <= "111111";
				when "1000000110001" => rgb <= "111111";
				when "1000000110010" => rgb <= "111111";
				when "1000000110011" => rgb <= "111111";
				when "1000000110100" => rgb <= "111111";
				when "1000000110101" => rgb <= "111111";
				when "1000000110110" => rgb <= "111111";
				when "1000000110111" => rgb <= "111111";
				when "1000010011000" => rgb <= "111111";
				when "1000010011001" => rgb <= "111111";
				when "1000010011010" => rgb <= "111111";
				when "1000010011011" => rgb <= "111111";
				when "1000010011100" => rgb <= "111111";
				when "1000010011101" => rgb <= "111111";
				when "1000010011110" => rgb <= "111111";
				when "1000010011111" => rgb <= "111111";
				when "1000010100000" => rgb <= "111111";
				when "1000010100001" => rgb <= "111111";
				when "1000010100010" => rgb <= "111111";
				when "1000010100011" => rgb <= "111111";
				when "1000010100100" => rgb <= "111111";
				when "1000010100101" => rgb <= "111111";
				when "1000010100110" => rgb <= "111111";
				when "1000010100111" => rgb <= "111111";
				when "1000010101000" => rgb <= "111111";
				when "1000010101001" => rgb <= "111111";
				when "1000010101010" => rgb <= "111111";
				when "1000010101011" => rgb <= "111111";
				when "1000010101100" => rgb <= "111111";
				when "1000010101101" => rgb <= "111111";
				when "1000010101110" => rgb <= "111111";
				when "1000010101111" => rgb <= "111111";
				when "1000010110000" => rgb <= "111111";
				when "1000010110001" => rgb <= "111111";
				when "1000010110010" => rgb <= "111111";
				when "1000010110011" => rgb <= "111111";
				when "1000010110100" => rgb <= "111111";
				when "1000010110101" => rgb <= "111111";
				when "1000010110110" => rgb <= "111111";
				when "1000010110111" => rgb <= "111111";
				when "1000100011000" => rgb <= "111111";
				when "1000100011001" => rgb <= "111111";
				when "1000100011010" => rgb <= "111111";
				when "1000100011011" => rgb <= "111111";
				when "1000100011100" => rgb <= "111111";
				when "1000100011101" => rgb <= "111111";
				when "1000100011110" => rgb <= "111111";
				when "1000100011111" => rgb <= "111111";
				when "1000100100000" => rgb <= "111111";
				when "1000100100001" => rgb <= "111111";
				when "1000100100010" => rgb <= "111111";
				when "1000100100011" => rgb <= "111111";
				when "1000100100100" => rgb <= "111111";
				when "1000100100101" => rgb <= "111111";
				when "1000100100110" => rgb <= "111111";
				when "1000100100111" => rgb <= "111111";
				when "1000100101000" => rgb <= "111111";
				when "1000100101001" => rgb <= "111111";
				when "1000100101010" => rgb <= "111111";
				when "1000100101011" => rgb <= "111111";
				when "1000100101100" => rgb <= "111111";
				when "1000100101101" => rgb <= "111111";
				when "1000100101110" => rgb <= "111111";
				when "1000100101111" => rgb <= "111111";
				when "1000100110000" => rgb <= "111111";
				when "1000100110001" => rgb <= "111111";
				when "1000100110010" => rgb <= "111111";
				when "1000100110011" => rgb <= "111111";
				when "1000100110100" => rgb <= "111111";
				when "1000100110101" => rgb <= "111111";
				when "1000100110110" => rgb <= "111111";
				when "1000100110111" => rgb <= "111111";
				when "1000110011000" => rgb <= "111111";
				when "1000110011001" => rgb <= "111111";
				when "1000110011010" => rgb <= "111111";
				when "1000110011011" => rgb <= "111111";
				when "1000110011100" => rgb <= "111111";
				when "1000110011101" => rgb <= "111111";
				when "1000110011110" => rgb <= "111111";
				when "1000110011111" => rgb <= "111111";
				when "1000110100000" => rgb <= "111111";
				when "1000110100001" => rgb <= "111111";
				when "1000110100010" => rgb <= "111111";
				when "1000110100011" => rgb <= "111111";
				when "1000110100100" => rgb <= "111111";
				when "1000110100101" => rgb <= "111111";
				when "1000110100110" => rgb <= "111111";
				when "1000110100111" => rgb <= "111111";
				when "1000110101000" => rgb <= "111111";
				when "1000110101001" => rgb <= "111111";
				when "1000110101010" => rgb <= "111111";
				when "1000110101011" => rgb <= "111111";
				when "1000110101100" => rgb <= "111111";
				when "1000110101101" => rgb <= "111111";
				when "1000110101110" => rgb <= "111111";
				when "1000110101111" => rgb <= "111111";
				when "1000110110000" => rgb <= "111111";
				when "1000110110001" => rgb <= "111111";
				when "1000110110010" => rgb <= "111111";
				when "1000110110011" => rgb <= "111111";
				when "1000110110100" => rgb <= "111111";
				when "1000110110101" => rgb <= "111111";
				when "1000110110110" => rgb <= "111111";
				when "1000110110111" => rgb <= "111111";
				when "1001000011000" => rgb <= "111111";
				when "1001000011001" => rgb <= "111111";
				when "1001000011100" => rgb <= "111111";
				when "1001000011101" => rgb <= "111111";
				when "1001000100000" => rgb <= "111111";
				when "1001000100001" => rgb <= "111111";
				when "1001000100100" => rgb <= "111111";
				when "1001000100101" => rgb <= "111111";
				when "1001000100110" => rgb <= "111111";
				when "1001000101001" => rgb <= "111111";
				when "1001000101010" => rgb <= "111111";
				when "1001000101011" => rgb <= "111111";
				when "1001000101110" => rgb <= "111111";
				when "1001000101111" => rgb <= "111111";
				when "1001000110010" => rgb <= "111111";
				when "1001000110011" => rgb <= "111111";
				when "1001000110110" => rgb <= "111111";
				when "1001000110111" => rgb <= "111111";
				when "1001010011000" => rgb <= "111111";
				when "1001010011001" => rgb <= "111111";
				when "1001010011100" => rgb <= "111111";
				when "1001010011101" => rgb <= "111111";
				when "1001010100000" => rgb <= "111111";
				when "1001010100001" => rgb <= "111111";
				when "1001010100100" => rgb <= "111111";
				when "1001010100101" => rgb <= "111111";
				when "1001010100110" => rgb <= "111111";
				when "1001010101001" => rgb <= "111111";
				when "1001010101010" => rgb <= "111111";
				when "1001010101011" => rgb <= "111111";
				when "1001010101110" => rgb <= "111111";
				when "1001010101111" => rgb <= "111111";
				when "1001010110010" => rgb <= "111111";
				when "1001010110011" => rgb <= "111111";
				when "1001010110110" => rgb <= "111111";
				when "1001010110111" => rgb <= "111111";
				when "1001100011000" => rgb <= "111111";
				when "1001100011001" => rgb <= "111111";
				when "1001100011100" => rgb <= "111111";
				when "1001100011101" => rgb <= "111111";
				when "1001100100000" => rgb <= "111111";
				when "1001100100001" => rgb <= "111111";
				when "1001100100100" => rgb <= "111111";
				when "1001100100101" => rgb <= "111111";
				when "1001100100110" => rgb <= "111111";
				when "1001100101001" => rgb <= "111111";
				when "1001100101010" => rgb <= "111111";
				when "1001100101011" => rgb <= "111111";
				when "1001100101110" => rgb <= "111111";
				when "1001100101111" => rgb <= "111111";
				when "1001100110010" => rgb <= "111111";
				when "1001100110011" => rgb <= "111111";
				when "1001100110110" => rgb <= "111111";
				when "1001100110111" => rgb <= "111111";
				when "1001110011000" => rgb <= "111111";
				when "1001110011001" => rgb <= "111111";
				when "1001110011100" => rgb <= "111111";
				when "1001110011101" => rgb <= "111111";
				when "1001110100000" => rgb <= "111111";
				when "1001110100001" => rgb <= "111111";
				when "1001110100100" => rgb <= "111111";
				when "1001110100101" => rgb <= "111111";
				when "1001110100110" => rgb <= "111111";
				when "1001110101001" => rgb <= "111111";
				when "1001110101010" => rgb <= "111111";
				when "1001110101011" => rgb <= "111111";
				when "1001110101110" => rgb <= "111111";
				when "1001110101111" => rgb <= "111111";
				when "1001110110010" => rgb <= "111111";
				when "1001110110011" => rgb <= "111111";
				when "1001110110110" => rgb <= "111111";
				when "1001110110111" => rgb <= "111111";
				when "1010000011000" => rgb <= "111111";
				when "1010000011001" => rgb <= "111111";
				when "1010000011100" => rgb <= "111111";
				when "1010000011101" => rgb <= "111111";
				when "1010000100000" => rgb <= "111111";
				when "1010000100001" => rgb <= "111111";
				when "1010000100100" => rgb <= "111111";
				when "1010000100101" => rgb <= "111111";
				when "1010000100110" => rgb <= "111111";
				when "1010000101001" => rgb <= "111111";
				when "1010000101010" => rgb <= "111111";
				when "1010000101011" => rgb <= "111111";
				when "1010000101110" => rgb <= "111111";
				when "1010000101111" => rgb <= "111111";
				when "1010000110010" => rgb <= "111111";
				when "1010000110011" => rgb <= "111111";
				when "1010000110110" => rgb <= "111111";
				when "1010000110111" => rgb <= "111111";
				when "1010010011000" => rgb <= "111111";
				when "1010010011001" => rgb <= "111111";
				when "1010010011100" => rgb <= "111111";
				when "1010010011101" => rgb <= "111111";
				when "1010010100000" => rgb <= "111111";
				when "1010010100001" => rgb <= "111111";
				when "1010010100100" => rgb <= "111111";
				when "1010010100101" => rgb <= "111111";
				when "1010010100110" => rgb <= "111111";
				when "1010010101001" => rgb <= "111111";
				when "1010010101010" => rgb <= "111111";
				when "1010010101011" => rgb <= "111111";
				when "1010010101110" => rgb <= "111111";
				when "1010010101111" => rgb <= "111111";
				when "1010010110010" => rgb <= "111111";
				when "1010010110011" => rgb <= "111111";
				when "1010010110110" => rgb <= "111111";
				when "1010010110111" => rgb <= "111111";
				when "1010100011000" => rgb <= "111111";
				when "1010100011001" => rgb <= "111111";
				when "1010100011010" => rgb <= "111111";
				when "1010100011011" => rgb <= "111111";
				when "1010100011100" => rgb <= "111111";
				when "1010100011101" => rgb <= "111111";
				when "1010100011110" => rgb <= "111111";
				when "1010100011111" => rgb <= "111111";
				when "1010100100000" => rgb <= "111111";
				when "1010100100001" => rgb <= "111111";
				when "1010100100010" => rgb <= "111111";
				when "1010100100011" => rgb <= "111111";
				when "1010100100100" => rgb <= "111111";
				when "1010100100101" => rgb <= "111111";
				when "1010100100110" => rgb <= "111111";
				when "1010100100111" => rgb <= "111111";
				when "1010100101000" => rgb <= "111111";
				when "1010100101001" => rgb <= "111111";
				when "1010100101010" => rgb <= "111111";
				when "1010100101011" => rgb <= "111111";
				when "1010100101100" => rgb <= "111111";
				when "1010100101101" => rgb <= "111111";
				when "1010100101110" => rgb <= "111111";
				when "1010100101111" => rgb <= "111111";
				when "1010100110000" => rgb <= "111111";
				when "1010100110001" => rgb <= "111111";
				when "1010100110010" => rgb <= "111111";
				when "1010100110011" => rgb <= "111111";
				when "1010100110100" => rgb <= "111111";
				when "1010100110101" => rgb <= "111111";
				when "1010100110110" => rgb <= "111111";
				when "1010100110111" => rgb <= "111111";
				when "1010110011000" => rgb <= "111111";
				when "1010110011001" => rgb <= "111111";
				when "1010110011010" => rgb <= "111111";
				when "1010110011011" => rgb <= "111111";
				when "1010110011100" => rgb <= "111111";
				when "1010110011101" => rgb <= "111111";
				when "1010110011110" => rgb <= "111111";
				when "1010110011111" => rgb <= "111111";
				when "1010110100000" => rgb <= "111111";
				when "1010110100001" => rgb <= "111111";
				when "1010110100010" => rgb <= "111111";
				when "1010110100011" => rgb <= "111111";
				when "1010110100100" => rgb <= "111111";
				when "1010110100101" => rgb <= "111111";
				when "1010110100110" => rgb <= "111111";
				when "1010110100111" => rgb <= "111111";
				when "1010110101000" => rgb <= "111111";
				when "1010110101001" => rgb <= "111111";
				when "1010110101010" => rgb <= "111111";
				when "1010110101011" => rgb <= "111111";
				when "1010110101100" => rgb <= "111111";
				when "1010110101101" => rgb <= "111111";
				when "1010110101110" => rgb <= "111111";
				when "1010110101111" => rgb <= "111111";
				when "1010110110000" => rgb <= "111111";
				when "1010110110001" => rgb <= "111111";
				when "1010110110010" => rgb <= "111111";
				when "1010110110011" => rgb <= "111111";
				when "1010110110100" => rgb <= "111111";
				when "1010110110101" => rgb <= "111111";
				when "1010110110110" => rgb <= "111111";
				when "1010110110111" => rgb <= "111111";
				when "1011000011000" => rgb <= "111111";
				when "1011000011001" => rgb <= "111111";
				when "1011000011010" => rgb <= "111111";
				when "1011000011011" => rgb <= "111111";
				when "1011000011100" => rgb <= "111111";
				when "1011000011101" => rgb <= "111111";
				when "1011000011110" => rgb <= "111111";
				when "1011000011111" => rgb <= "111111";
				when "1011000100000" => rgb <= "111111";
				when "1011000100001" => rgb <= "111111";
				when "1011000100010" => rgb <= "111111";
				when "1011000100011" => rgb <= "111111";
				when "1011000100100" => rgb <= "111111";
				when "1011000100101" => rgb <= "111111";
				when "1011000100110" => rgb <= "111111";
				when "1011000100111" => rgb <= "111111";
				when "1011000101000" => rgb <= "111111";
				when "1011000101001" => rgb <= "111111";
				when "1011000101010" => rgb <= "111111";
				when "1011000101011" => rgb <= "111111";
				when "1011000101100" => rgb <= "111111";
				when "1011000101101" => rgb <= "111111";
				when "1011000101110" => rgb <= "111111";
				when "1011000101111" => rgb <= "111111";
				when "1011000110000" => rgb <= "111111";
				when "1011000110001" => rgb <= "111111";
				when "1011000110010" => rgb <= "111111";
				when "1011000110011" => rgb <= "111111";
				when "1011000110100" => rgb <= "111111";
				when "1011000110101" => rgb <= "111111";
				when "1011000110110" => rgb <= "111111";
				when "1011000110111" => rgb <= "111111";
				when "1011010011000" => rgb <= "111111";
				when "1011010011001" => rgb <= "111111";
				when "1011010011010" => rgb <= "111111";
				when "1011010011011" => rgb <= "111111";
				when "1011010011100" => rgb <= "111111";
				when "1011010011101" => rgb <= "111111";
				when "1011010011110" => rgb <= "111111";
				when "1011010011111" => rgb <= "111111";
				when "1011010100000" => rgb <= "111111";
				when "1011010100001" => rgb <= "111111";
				when "1011010100010" => rgb <= "111111";
				when "1011010100011" => rgb <= "111111";
				when "1011010100100" => rgb <= "111111";
				when "1011010100101" => rgb <= "111111";
				when "1011010100110" => rgb <= "111111";
				when "1011010100111" => rgb <= "111111";
				when "1011010101000" => rgb <= "111111";
				when "1011010101001" => rgb <= "111111";
				when "1011010101010" => rgb <= "111111";
				when "1011010101011" => rgb <= "111111";
				when "1011010101100" => rgb <= "111111";
				when "1011010101101" => rgb <= "111111";
				when "1011010101110" => rgb <= "111111";
				when "1011010101111" => rgb <= "111111";
				when "1011010110000" => rgb <= "111111";
				when "1011010110001" => rgb <= "111111";
				when "1011010110010" => rgb <= "111111";
				when "1011010110011" => rgb <= "111111";
				when "1011010110100" => rgb <= "111111";
				when "1011010110101" => rgb <= "111111";
				when "1011010110110" => rgb <= "111111";
				when "1011010110111" => rgb <= "111111";
				when "1011100011000" => rgb <= "111111";
				when "1011100011001" => rgb <= "111111";
				when "1011100011110" => rgb <= "111111";
				when "1011100011111" => rgb <= "111111";
				when "1011100100000" => rgb <= "111111";
				when "1011100100001" => rgb <= "111111";
				when "1011100100010" => rgb <= "111111";
				when "1011100100011" => rgb <= "111111";
				when "1011100100100" => rgb <= "111111";
				when "1011100100101" => rgb <= "111111";
				when "1011100101010" => rgb <= "111111";
				when "1011100101011" => rgb <= "111111";
				when "1011100110000" => rgb <= "111111";
				when "1011100110001" => rgb <= "111111";
				when "1011100110110" => rgb <= "111111";
				when "1011100110111" => rgb <= "111111";
				when "1011110000100" => rgb <= "111111";
				when "1011110000101" => rgb <= "111111";
				when "1011110000110" => rgb <= "111111";
				when "1011110000111" => rgb <= "111111";
				when "1011110001000" => rgb <= "111111";
				when "1011110011000" => rgb <= "111111";
				when "1011110011001" => rgb <= "111111";
				when "1011110011110" => rgb <= "111111";
				when "1011110011111" => rgb <= "111111";
				when "1011110100000" => rgb <= "111111";
				when "1011110100001" => rgb <= "111111";
				when "1011110100010" => rgb <= "111111";
				when "1011110100011" => rgb <= "111111";
				when "1011110100100" => rgb <= "111111";
				when "1011110100101" => rgb <= "111111";
				when "1011110101010" => rgb <= "111111";
				when "1011110101011" => rgb <= "111111";
				when "1011110110000" => rgb <= "111111";
				when "1011110110001" => rgb <= "111111";
				when "1011110110110" => rgb <= "111111";
				when "1011110110111" => rgb <= "111111";
				when "1011111000111" => rgb <= "111111";
				when "1011111001000" => rgb <= "111111";
				when "1011111001001" => rgb <= "111111";
				when "1011111001010" => rgb <= "111111";
				when "1011111001011" => rgb <= "111111";
				when "1100000000011" => rgb <= "111111";
				when "1100000000100" => rgb <= "111111";
				when "1100000000101" => rgb <= "111111";
				when "1100000000110" => rgb <= "111111";
				when "1100000001000" => rgb <= "111111";
				when "1100000011000" => rgb <= "111111";
				when "1100000011001" => rgb <= "111111";
				when "1100000011110" => rgb <= "111111";
				when "1100000011111" => rgb <= "111111";
				when "1100000100000" => rgb <= "111111";
				when "1100000100001" => rgb <= "111111";
				when "1100000100010" => rgb <= "001011";
				when "1100000100011" => rgb <= "001011";
				when "1100000100100" => rgb <= "111111";
				when "1100000100101" => rgb <= "111111";
				when "1100000100110" => rgb <= "111111";
				when "1100000100111" => rgb <= "111111";
				when "1100000101000" => rgb <= "111111";
				when "1100000101001" => rgb <= "111111";
				when "1100000101010" => rgb <= "111111";
				when "1100000101011" => rgb <= "111111";
				when "1100000101100" => rgb <= "111111";
				when "1100000101101" => rgb <= "111111";
				when "1100000101110" => rgb <= "111111";
				when "1100000101111" => rgb <= "111111";
				when "1100000110000" => rgb <= "111111";
				when "1100000110001" => rgb <= "111111";
				when "1100000110010" => rgb <= "111111";
				when "1100000110011" => rgb <= "111111";
				when "1100000110100" => rgb <= "111111";
				when "1100000110101" => rgb <= "111111";
				when "1100000110110" => rgb <= "111111";
				when "1100000110111" => rgb <= "111111";
				when "1100001000111" => rgb <= "111111";
				when "1100001001001" => rgb <= "111111";
				when "1100001001010" => rgb <= "111111";
				when "1100001001011" => rgb <= "111111";
				when "1100001001100" => rgb <= "111111";
				when "1100010000010" => rgb <= "111111";
				when "1100010000011" => rgb <= "111111";
				when "1100010000100" => rgb <= "111111";
				when "1100010000101" => rgb <= "111111";
				when "1100010000110" => rgb <= "111111";
				when "1100010000111" => rgb <= "111111";
				when "1100010001000" => rgb <= "111111";
				when "1100010011000" => rgb <= "111111";
				when "1100010011001" => rgb <= "111111";
				when "1100010011110" => rgb <= "111111";
				when "1100010011111" => rgb <= "111111";
				when "1100010100000" => rgb <= "111111";
				when "1100010100001" => rgb <= "111111";
				when "1100010100010" => rgb <= "001011";
				when "1100010100011" => rgb <= "001011";
				when "1100010100100" => rgb <= "111111";
				when "1100010100101" => rgb <= "111111";
				when "1100010100110" => rgb <= "111111";
				when "1100010100111" => rgb <= "111111";
				when "1100010101000" => rgb <= "111111";
				when "1100010101001" => rgb <= "111111";
				when "1100010101010" => rgb <= "111111";
				when "1100010101011" => rgb <= "111111";
				when "1100010101100" => rgb <= "111111";
				when "1100010101101" => rgb <= "111111";
				when "1100010101110" => rgb <= "111111";
				when "1100010101111" => rgb <= "111111";
				when "1100010110000" => rgb <= "111111";
				when "1100010110001" => rgb <= "111111";
				when "1100010110010" => rgb <= "111111";
				when "1100010110011" => rgb <= "111111";
				when "1100010110100" => rgb <= "111111";
				when "1100010110101" => rgb <= "111111";
				when "1100010110110" => rgb <= "111111";
				when "1100010110111" => rgb <= "111111";
				when "1100011000111" => rgb <= "111111";
				when "1100011001000" => rgb <= "111111";
				when "1100011001001" => rgb <= "111111";
				when "1100011001010" => rgb <= "111111";
				when "1100011001011" => rgb <= "111111";
				when "1100011001100" => rgb <= "111111";
				when "1100011001101" => rgb <= "111111";
				when "1100100000011" => rgb <= "111111";
				when "1100100000100" => rgb <= "111111";
				when "1100100000101" => rgb <= "111111";
				when "1100100000110" => rgb <= "111111";
				when "1100100000111" => rgb <= "111111";
				when "1100100001000" => rgb <= "111111";
				when "1100100011000" => rgb <= "111111";
				when "1100100011001" => rgb <= "111111";
				when "1100100011010" => rgb <= "111111";
				when "1100100011011" => rgb <= "111111";
				when "1100100011100" => rgb <= "111111";
				when "1100100011101" => rgb <= "111111";
				when "1100100011110" => rgb <= "111111";
				when "1100100011111" => rgb <= "111111";
				when "1100100100000" => rgb <= "111111";
				when "1100100100001" => rgb <= "111111";
				when "1100100100010" => rgb <= "001011";
				when "1100100100011" => rgb <= "001011";
				when "1100100100100" => rgb <= "111111";
				when "1100100100101" => rgb <= "111111";
				when "1100100100110" => rgb <= "111111";
				when "1100100100111" => rgb <= "111111";
				when "1100100101000" => rgb <= "111111";
				when "1100100101001" => rgb <= "111111";
				when "1100100101010" => rgb <= "111111";
				when "1100100101011" => rgb <= "111111";
				when "1100100101100" => rgb <= "111111";
				when "1100100101101" => rgb <= "111111";
				when "1100100101110" => rgb <= "111111";
				when "1100100101111" => rgb <= "111111";
				when "1100100110000" => rgb <= "111111";
				when "1100100110001" => rgb <= "111111";
				when "1100100110010" => rgb <= "111111";
				when "1100100110011" => rgb <= "111111";
				when "1100100110100" => rgb <= "111111";
				when "1100100110101" => rgb <= "111111";
				when "1100100110110" => rgb <= "111111";
				when "1100100110111" => rgb <= "111111";
				when "1100101000111" => rgb <= "111111";
				when "1100101001000" => rgb <= "111111";
				when "1100101001001" => rgb <= "111111";
				when "1100101001010" => rgb <= "111111";
				when "1100101001011" => rgb <= "111111";
				when "1100101001100" => rgb <= "111111";
				when "1100110000011" => rgb <= "111111";
				when "1100110000100" => rgb <= "111111";
				when "1100110000110" => rgb <= "111111";
				when "1100110000111" => rgb <= "111111";
				when "1100110011000" => rgb <= "111111";
				when "1100110011001" => rgb <= "111111";
				when "1100110011010" => rgb <= "111111";
				when "1100110011011" => rgb <= "111111";
				when "1100110011100" => rgb <= "111111";
				when "1100110011101" => rgb <= "111111";
				when "1100110011110" => rgb <= "111111";
				when "1100110011111" => rgb <= "111111";
				when "1100110100000" => rgb <= "111111";
				when "1100110100001" => rgb <= "111111";
				when "1100110100010" => rgb <= "001011";
				when "1100110100011" => rgb <= "001011";
				when "1100110100100" => rgb <= "111111";
				when "1100110100101" => rgb <= "111111";
				when "1100110100110" => rgb <= "111111";
				when "1100110100111" => rgb <= "111111";
				when "1100110101000" => rgb <= "111111";
				when "1100110101001" => rgb <= "111111";
				when "1100110101010" => rgb <= "111111";
				when "1100110101011" => rgb <= "111111";
				when "1100110101100" => rgb <= "111111";
				when "1100110101101" => rgb <= "111111";
				when "1100110101110" => rgb <= "111111";
				when "1100110101111" => rgb <= "111111";
				when "1100110110000" => rgb <= "111111";
				when "1100110110001" => rgb <= "111111";
				when "1100110110010" => rgb <= "111111";
				when "1100110110011" => rgb <= "111111";
				when "1100110110100" => rgb <= "111111";
				when "1100110110101" => rgb <= "111111";
				when "1100110110110" => rgb <= "111111";
				when "1100110110111" => rgb <= "111111";
				when "1100111001000" => rgb <= "111111";
				when "1100111001001" => rgb <= "111111";
				when "1100111001011" => rgb <= "111111";
				when "1100111001100" => rgb <= "111111";
				when "1101000000000" => rgb <= "111111";
				when "1101000000001" => rgb <= "111111";
				when "1101000000010" => rgb <= "111111";
				when "1101000000011" => rgb <= "111111";
				when "1101000000100" => rgb <= "111111";
				when "1101000000101" => rgb <= "111111";
				when "1101000000110" => rgb <= "111111";
				when "1101000000111" => rgb <= "111111";
				when "1101000001000" => rgb <= "111111";
				when "1101000001001" => rgb <= "111111";
				when "1101000001010" => rgb <= "111111";
				when "1101000001011" => rgb <= "111111";
				when "1101000001100" => rgb <= "111111";
				when "1101000001101" => rgb <= "111111";
				when "1101000001110" => rgb <= "111111";
				when "1101000001111" => rgb <= "111111";
				when "1101000010000" => rgb <= "111111";
				when "1101000010001" => rgb <= "111111";
				when "1101000010010" => rgb <= "111111";
				when "1101000010011" => rgb <= "111111";
				when "1101000010100" => rgb <= "111111";
				when "1101000010101" => rgb <= "111111";
				when "1101000010110" => rgb <= "111111";
				when "1101000010111" => rgb <= "111111";
				when "1101000011000" => rgb <= "111111";
				when "1101000011001" => rgb <= "111111";
				when "1101000011010" => rgb <= "111111";
				when "1101000011011" => rgb <= "111111";
				when "1101000011100" => rgb <= "111111";
				when "1101000011101" => rgb <= "111111";
				when "1101000011110" => rgb <= "111111";
				when "1101000011111" => rgb <= "111111";
				when "1101000100000" => rgb <= "111111";
				when "1101000100001" => rgb <= "111111";
				when "1101000100010" => rgb <= "111111";
				when "1101000100011" => rgb <= "111111";
				when "1101000100100" => rgb <= "111111";
				when "1101000100101" => rgb <= "111111";
				when "1101000100110" => rgb <= "111111";
				when "1101000100111" => rgb <= "111111";
				when "1101000101000" => rgb <= "111111";
				when "1101000101001" => rgb <= "111111";
				when "1101000101010" => rgb <= "111111";
				when "1101000101011" => rgb <= "111111";
				when "1101000101100" => rgb <= "111111";
				when "1101000101101" => rgb <= "111111";
				when "1101000101110" => rgb <= "111111";
				when "1101000101111" => rgb <= "111111";
				when "1101000110000" => rgb <= "111111";
				when "1101000110001" => rgb <= "111111";
				when "1101000110010" => rgb <= "111111";
				when "1101000110011" => rgb <= "111111";
				when "1101000110100" => rgb <= "111111";
				when "1101000110101" => rgb <= "111111";
				when "1101000110110" => rgb <= "111111";
				when "1101000110111" => rgb <= "111111";
				when "1101000111000" => rgb <= "111111";
				when "1101000111001" => rgb <= "111111";
				when "1101000111010" => rgb <= "111111";
				when "1101000111011" => rgb <= "111111";
				when "1101000111100" => rgb <= "111111";
				when "1101000111101" => rgb <= "111111";
				when "1101000111110" => rgb <= "111111";
				when "1101000111111" => rgb <= "111111";
				when "1101001000000" => rgb <= "111111";
				when "1101001000001" => rgb <= "111111";
				when "1101001000010" => rgb <= "111111";
				when "1101001000011" => rgb <= "111111";
				when "1101001000100" => rgb <= "111111";
				when "1101001000101" => rgb <= "111111";
				when "1101001000110" => rgb <= "111111";
				when "1101001000111" => rgb <= "111111";
				when "1101001001000" => rgb <= "111111";
				when "1101001001001" => rgb <= "111111";
				when "1101001001010" => rgb <= "111111";
				when "1101001001011" => rgb <= "111111";
				when "1101001001100" => rgb <= "111111";
				when "1101001001101" => rgb <= "111111";
				when "1101001001110" => rgb <= "111111";
				when "1101001001111" => rgb <= "111111";
				when "1101010000000" => rgb <= "111111";
				when "1101010000001" => rgb <= "111111";
				when "1101010000010" => rgb <= "111111";
				when "1101010000011" => rgb <= "111111";
				when "1101010000100" => rgb <= "111111";
				when "1101010000101" => rgb <= "111111";
				when "1101010000110" => rgb <= "111111";
				when "1101010000111" => rgb <= "111111";
				when "1101010001000" => rgb <= "111111";
				when "1101010001001" => rgb <= "111111";
				when "1101010001010" => rgb <= "111111";
				when "1101010001011" => rgb <= "111111";
				when "1101010001100" => rgb <= "111111";
				when "1101010001101" => rgb <= "111111";
				when "1101010001110" => rgb <= "111111";
				when "1101010001111" => rgb <= "111111";
				when "1101010010000" => rgb <= "111111";
				when "1101010010001" => rgb <= "111111";
				when "1101010010010" => rgb <= "111111";
				when "1101010010011" => rgb <= "111111";
				when "1101010010100" => rgb <= "111111";
				when "1101010010101" => rgb <= "111111";
				when "1101010010110" => rgb <= "111111";
				when "1101010010111" => rgb <= "111111";
				when "1101010011000" => rgb <= "111111";
				when "1101010011001" => rgb <= "111111";
				when "1101010011010" => rgb <= "111111";
				when "1101010011011" => rgb <= "111111";
				when "1101010011100" => rgb <= "111111";
				when "1101010011101" => rgb <= "111111";
				when "1101010011110" => rgb <= "111111";
				when "1101010011111" => rgb <= "111111";
				when "1101010100000" => rgb <= "111111";
				when "1101010100001" => rgb <= "111111";
				when "1101010100010" => rgb <= "111111";
				when "1101010100011" => rgb <= "111111";
				when "1101010100100" => rgb <= "111111";
				when "1101010100101" => rgb <= "111111";
				when "1101010100110" => rgb <= "111111";
				when "1101010100111" => rgb <= "111111";
				when "1101010101000" => rgb <= "111111";
				when "1101010101001" => rgb <= "111111";
				when "1101010101010" => rgb <= "111111";
				when "1101010101011" => rgb <= "111111";
				when "1101010101100" => rgb <= "111111";
				when "1101010101101" => rgb <= "111111";
				when "1101010101110" => rgb <= "111111";
				when "1101010101111" => rgb <= "111111";
				when "1101010110000" => rgb <= "111111";
				when "1101010110001" => rgb <= "111111";
				when "1101010110010" => rgb <= "111111";
				when "1101010110011" => rgb <= "111111";
				when "1101010110100" => rgb <= "111111";
				when "1101010110101" => rgb <= "111111";
				when "1101010110110" => rgb <= "111111";
				when "1101010110111" => rgb <= "111111";
				when "1101010111000" => rgb <= "111111";
				when "1101010111001" => rgb <= "111111";
				when "1101010111010" => rgb <= "111111";
				when "1101010111011" => rgb <= "111111";
				when "1101010111100" => rgb <= "111111";
				when "1101010111101" => rgb <= "111111";
				when "1101010111110" => rgb <= "111111";
				when "1101010111111" => rgb <= "111111";
				when "1101011000000" => rgb <= "111111";
				when "1101011000001" => rgb <= "111111";
				when "1101011000010" => rgb <= "111111";
				when "1101011000011" => rgb <= "111111";
				when "1101011000100" => rgb <= "111111";
				when "1101011000101" => rgb <= "111111";
				when "1101011000110" => rgb <= "111111";
				when "1101011000111" => rgb <= "111111";
				when "1101011001000" => rgb <= "111111";
				when "1101011001001" => rgb <= "111111";
				when "1101011001010" => rgb <= "111111";
				when "1101011001011" => rgb <= "111111";
				when "1101011001100" => rgb <= "111111";
				when "1101011001101" => rgb <= "111111";
				when "1101011001110" => rgb <= "111111";
				when "1101011001111" => rgb <= "111111";
				when "1101110000000" => rgb <= "111000";
				when "1101110000001" => rgb <= "111000";
				when "1101110000010" => rgb <= "111000";
				when "1101110000011" => rgb <= "111000";
				when "1101110000100" => rgb <= "111000";
				when "1101110000101" => rgb <= "111000";
				when "1101110000110" => rgb <= "111000";
				when "1101110000111" => rgb <= "111000";
				when "1101110001000" => rgb <= "111000";
				when "1101110001001" => rgb <= "111000";
				when "1101110001010" => rgb <= "111000";
				when "1101110001011" => rgb <= "111000";
				when "1101110001100" => rgb <= "111000";
				when "1101110001101" => rgb <= "111000";
				when "1101110001110" => rgb <= "111000";
				when "1101110001111" => rgb <= "111000";
				when "1101110010000" => rgb <= "111000";
				when "1101110010001" => rgb <= "111000";
				when "1101110010010" => rgb <= "111000";
				when "1101110010011" => rgb <= "111000";
				when "1101110010100" => rgb <= "111000";
				when "1101110010101" => rgb <= "111000";
				when "1101110010110" => rgb <= "111000";
				when "1101110010111" => rgb <= "111000";
				when "1101110011000" => rgb <= "111000";
				when "1101110011001" => rgb <= "111000";
				when "1101110011010" => rgb <= "111000";
				when "1101110011011" => rgb <= "111000";
				when "1101110011100" => rgb <= "111000";
				when "1101110011101" => rgb <= "111000";
				when "1101110011110" => rgb <= "111000";
				when "1101110011111" => rgb <= "111000";
				when "1101110100000" => rgb <= "111000";
				when "1101110100001" => rgb <= "111000";
				when "1101110100010" => rgb <= "111000";
				when "1101110100011" => rgb <= "111000";
				when "1101110100100" => rgb <= "111000";
				when "1101110100101" => rgb <= "111000";
				when "1101110100110" => rgb <= "111000";
				when "1101110100111" => rgb <= "111000";
				when "1101110101000" => rgb <= "111000";
				when "1101110101001" => rgb <= "111000";
				when "1101110101010" => rgb <= "111000";
				when "1101110101011" => rgb <= "111000";
				when "1101110101100" => rgb <= "111000";
				when "1101110101101" => rgb <= "111000";
				when "1101110101110" => rgb <= "111000";
				when "1101110101111" => rgb <= "111000";
				when "1101110110000" => rgb <= "111000";
				when "1101110110001" => rgb <= "111000";
				when "1101110110010" => rgb <= "111000";
				when "1101110110011" => rgb <= "111000";
				when "1101110110100" => rgb <= "111000";
				when "1101110110101" => rgb <= "111000";
				when "1101110110110" => rgb <= "111000";
				when "1101110110111" => rgb <= "111000";
				when "1101110111000" => rgb <= "111000";
				when "1101110111001" => rgb <= "111000";
				when "1101110111010" => rgb <= "111000";
				when "1101110111011" => rgb <= "111000";
				when "1101110111100" => rgb <= "111000";
				when "1101110111101" => rgb <= "111000";
				when "1101110111110" => rgb <= "111000";
				when "1101110111111" => rgb <= "111000";
				when "1101111000000" => rgb <= "111000";
				when "1101111000001" => rgb <= "111000";
				when "1101111000010" => rgb <= "111000";
				when "1101111000011" => rgb <= "111000";
				when "1101111000100" => rgb <= "111000";
				when "1101111000101" => rgb <= "111000";
				when "1101111000110" => rgb <= "111000";
				when "1101111000111" => rgb <= "111000";
				when "1101111001000" => rgb <= "111000";
				when "1101111001001" => rgb <= "111000";
				when "1101111001010" => rgb <= "111000";
				when "1101111001011" => rgb <= "111000";
				when "1101111001100" => rgb <= "111000";
				when "1101111001101" => rgb <= "111000";
				when "1101111001110" => rgb <= "111000";
				when "1101111001111" => rgb <= "111000";
				when "1110010000000" => rgb <= "111111";
				when "1110010000001" => rgb <= "111111";
				when "1110010000010" => rgb <= "111111";
				when "1110010000011" => rgb <= "111111";
				when "1110010000100" => rgb <= "111111";
				when "1110010000101" => rgb <= "111111";
				when "1110010000110" => rgb <= "111111";
				when "1110010000111" => rgb <= "111111";
				when "1110010001000" => rgb <= "111111";
				when "1110010001001" => rgb <= "111111";
				when "1110010001010" => rgb <= "111111";
				when "1110010001011" => rgb <= "111111";
				when "1110010001100" => rgb <= "111111";
				when "1110010001101" => rgb <= "111111";
				when "1110010001110" => rgb <= "111111";
				when "1110010001111" => rgb <= "111111";
				when "1110010010000" => rgb <= "111111";
				when "1110010010001" => rgb <= "111111";
				when "1110010010010" => rgb <= "111111";
				when "1110010010011" => rgb <= "111111";
				when "1110010010100" => rgb <= "111111";
				when "1110010010101" => rgb <= "111111";
				when "1110010010110" => rgb <= "111111";
				when "1110010010111" => rgb <= "111111";
				when "1110010011000" => rgb <= "111111";
				when "1110010011001" => rgb <= "111111";
				when "1110010011010" => rgb <= "111111";
				when "1110010011011" => rgb <= "111111";
				when "1110010011100" => rgb <= "111111";
				when "1110010011101" => rgb <= "111111";
				when "1110010011110" => rgb <= "111111";
				when "1110010011111" => rgb <= "111111";
				when "1110010100000" => rgb <= "111111";
				when "1110010100001" => rgb <= "111111";
				when "1110010100010" => rgb <= "111111";
				when "1110010100011" => rgb <= "111111";
				when "1110010100100" => rgb <= "111111";
				when "1110010100101" => rgb <= "111111";
				when "1110010100110" => rgb <= "111111";
				when "1110010100111" => rgb <= "111111";
				when "1110010101000" => rgb <= "111111";
				when "1110010101001" => rgb <= "111111";
				when "1110010101010" => rgb <= "111111";
				when "1110010101011" => rgb <= "111111";
				when "1110010101100" => rgb <= "111111";
				when "1110010101101" => rgb <= "111111";
				when "1110010101110" => rgb <= "111111";
				when "1110010101111" => rgb <= "111111";
				when "1110010110000" => rgb <= "111111";
				when "1110010110001" => rgb <= "111111";
				when "1110010110010" => rgb <= "111111";
				when "1110010110011" => rgb <= "111111";
				when "1110010110100" => rgb <= "111111";
				when "1110010110101" => rgb <= "111111";
				when "1110010110110" => rgb <= "111111";
				when "1110010110111" => rgb <= "111111";
				when "1110010111000" => rgb <= "111111";
				when "1110010111001" => rgb <= "111111";
				when "1110010111010" => rgb <= "111111";
				when "1110010111011" => rgb <= "111111";
				when "1110010111100" => rgb <= "111111";
				when "1110010111101" => rgb <= "111111";
				when "1110010111110" => rgb <= "111111";
				when "1110010111111" => rgb <= "111111";
				when "1110011000000" => rgb <= "111111";
				when "1110011000001" => rgb <= "111111";
				when "1110011000010" => rgb <= "111111";
				when "1110011000011" => rgb <= "111111";
				when "1110011000100" => rgb <= "111111";
				when "1110011000101" => rgb <= "111111";
				when "1110011000110" => rgb <= "111111";
				when "1110011000111" => rgb <= "111111";
				when "1110011001000" => rgb <= "111111";
				when "1110011001001" => rgb <= "111111";
				when "1110011001010" => rgb <= "111111";
				when "1110011001011" => rgb <= "111111";
				when "1110011001100" => rgb <= "111111";
				when "1110011001101" => rgb <= "111111";
				when "1110011001110" => rgb <= "111111";
				when "1110011001111" => rgb <= "111111";
				when "1110100000000" => rgb <= "111111";
				when "1110100000001" => rgb <= "111111";
				when "1110100000010" => rgb <= "111111";
				when "1110100000011" => rgb <= "111111";
				when "1110100000100" => rgb <= "111111";
				when "1110100000101" => rgb <= "111111";
				when "1110100000110" => rgb <= "111111";
				when "1110100000111" => rgb <= "111111";
				when "1110100001000" => rgb <= "111111";
				when "1110100001001" => rgb <= "111111";
				when "1110100001010" => rgb <= "111111";
				when "1110100001011" => rgb <= "111111";
				when "1110100001100" => rgb <= "111111";
				when "1110100001101" => rgb <= "111111";
				when "1110100001110" => rgb <= "111111";
				when "1110100001111" => rgb <= "111111";
				when "1110100010000" => rgb <= "111111";
				when "1110100010001" => rgb <= "111111";
				when "1110100010010" => rgb <= "111111";
				when "1110100010011" => rgb <= "111111";
				when "1110100010100" => rgb <= "111111";
				when "1110100010101" => rgb <= "111111";
				when "1110100010110" => rgb <= "111111";
				when "1110100010111" => rgb <= "111111";
				when "1110100011000" => rgb <= "111111";
				when "1110100011001" => rgb <= "111111";
				when "1110100011010" => rgb <= "111111";
				when "1110100011011" => rgb <= "111111";
				when "1110100011100" => rgb <= "111111";
				when "1110100011101" => rgb <= "111111";
				when "1110100011110" => rgb <= "111111";
				when "1110100011111" => rgb <= "111111";
				when "1110100100000" => rgb <= "111111";
				when "1110100100001" => rgb <= "111111";
				when "1110100100010" => rgb <= "111111";
				when "1110100100011" => rgb <= "111111";
				when "1110100100100" => rgb <= "111111";
				when "1110100100101" => rgb <= "111111";
				when "1110100100110" => rgb <= "111111";
				when "1110100100111" => rgb <= "111111";
				when "1110100101000" => rgb <= "111111";
				when "1110100101001" => rgb <= "111111";
				when "1110100101010" => rgb <= "111111";
				when "1110100101011" => rgb <= "111111";
				when "1110100101100" => rgb <= "111111";
				when "1110100101101" => rgb <= "111111";
				when "1110100101110" => rgb <= "111111";
				when "1110100101111" => rgb <= "111111";
				when "1110100110000" => rgb <= "111111";
				when "1110100110001" => rgb <= "111111";
				when "1110100110010" => rgb <= "111111";
				when "1110100110011" => rgb <= "111111";
				when "1110100110100" => rgb <= "111111";
				when "1110100110101" => rgb <= "111111";
				when "1110100110110" => rgb <= "111111";
				when "1110100110111" => rgb <= "111111";
				when "1110100111000" => rgb <= "111111";
				when "1110100111001" => rgb <= "111111";
				when "1110100111010" => rgb <= "111111";
				when "1110100111011" => rgb <= "111111";
				when "1110100111100" => rgb <= "111111";
				when "1110100111101" => rgb <= "111111";
				when "1110100111110" => rgb <= "111111";
				when "1110100111111" => rgb <= "111111";
				when "1110101000000" => rgb <= "111111";
				when "1110101000001" => rgb <= "111111";
				when "1110101000010" => rgb <= "111111";
				when "1110101000011" => rgb <= "111111";
				when "1110101000100" => rgb <= "111111";
				when "1110101000101" => rgb <= "111111";
				when "1110101000110" => rgb <= "111111";
				when "1110101000111" => rgb <= "111111";
				when "1110101001000" => rgb <= "111111";
				when "1110101001001" => rgb <= "111111";
				when "1110101001010" => rgb <= "111111";
				when "1110101001011" => rgb <= "111111";
				when "1110101001100" => rgb <= "111111";
				when "1110101001101" => rgb <= "111111";
				when "1110101001110" => rgb <= "111111";
				when "1110101001111" => rgb <= "111111";
				when "1110110000000" => rgb <= "111111";
				when "1110110000001" => rgb <= "111111";
				when "1110110000010" => rgb <= "111111";
				when "1110110000011" => rgb <= "111111";
				when "1110110000100" => rgb <= "111111";
				when "1110110000101" => rgb <= "111111";
				when "1110110000110" => rgb <= "111111";
				when "1110110000111" => rgb <= "111111";
				when "1110110001000" => rgb <= "111111";
				when "1110110001001" => rgb <= "111111";
				when "1110110001010" => rgb <= "111111";
				when "1110110001011" => rgb <= "111111";
				when "1110110001100" => rgb <= "111111";
				when "1110110001101" => rgb <= "111111";
				when "1110110001110" => rgb <= "111111";
				when "1110110001111" => rgb <= "111111";
				when "1110110010000" => rgb <= "111111";
				when "1110110010001" => rgb <= "111111";
				when "1110110010010" => rgb <= "111111";
				when "1110110010011" => rgb <= "111111";
				when "1110110010100" => rgb <= "111111";
				when "1110110010101" => rgb <= "111111";
				when "1110110010110" => rgb <= "111111";
				when "1110110010111" => rgb <= "111111";
				when "1110110011000" => rgb <= "111111";
				when "1110110011001" => rgb <= "111111";
				when "1110110011010" => rgb <= "111111";
				when "1110110011011" => rgb <= "111111";
				when "1110110011100" => rgb <= "111111";
				when "1110110011101" => rgb <= "111111";
				when "1110110011110" => rgb <= "111111";
				when "1110110011111" => rgb <= "111111";
				when "1110110100000" => rgb <= "111111";
				when "1110110100001" => rgb <= "111111";
				when "1110110100010" => rgb <= "111111";
				when "1110110100011" => rgb <= "111111";
				when "1110110100100" => rgb <= "111111";
				when "1110110100101" => rgb <= "111111";
				when "1110110100110" => rgb <= "111111";
				when "1110110100111" => rgb <= "111111";
				when "1110110101000" => rgb <= "111111";
				when "1110110101001" => rgb <= "111111";
				when "1110110101010" => rgb <= "111111";
				when "1110110101011" => rgb <= "111111";
				when "1110110101100" => rgb <= "111111";
				when "1110110101101" => rgb <= "111111";
				when "1110110101110" => rgb <= "111111";
				when "1110110101111" => rgb <= "111111";
				when "1110110110000" => rgb <= "111111";
				when "1110110110001" => rgb <= "111111";
				when "1110110110010" => rgb <= "111111";
				when "1110110110011" => rgb <= "111111";
				when "1110110110100" => rgb <= "111111";
				when "1110110110101" => rgb <= "111111";
				when "1110110110110" => rgb <= "111111";
				when "1110110110111" => rgb <= "111111";
				when "1110110111000" => rgb <= "111111";
				when "1110110111001" => rgb <= "111111";
				when "1110110111010" => rgb <= "111111";
				when "1110110111011" => rgb <= "111111";
				when "1110110111100" => rgb <= "111111";
				when "1110110111101" => rgb <= "111111";
				when "1110110111110" => rgb <= "111111";
				when "1110110111111" => rgb <= "111111";
				when "1110111000000" => rgb <= "111111";
				when "1110111000001" => rgb <= "111111";
				when "1110111000010" => rgb <= "111111";
				when "1110111000011" => rgb <= "111111";
				when "1110111000100" => rgb <= "111111";
				when "1110111000101" => rgb <= "111111";
				when "1110111000110" => rgb <= "111111";
				when "1110111000111" => rgb <= "111111";
				when "1110111001000" => rgb <= "111111";
				when "1110111001001" => rgb <= "111111";
				when "1110111001010" => rgb <= "111111";
				when "1110111001011" => rgb <= "111111";
				when "1110111001100" => rgb <= "111111";
				when "1110111001101" => rgb <= "111111";
				when "1110111001110" => rgb <= "111111";
				when "1110111001111" => rgb <= "111111";
				when others => rgb <= "000000";
			end case;
		end if;
	end process;
	location <= std_logic_vector(col_idx) & std_logic_vector(row_idx);
end;
