library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity background_rom is
  port(
	  clk : in std_logic;
	  row_idx: in unsigned(7 downto 0);
	  col_idx : in unsigned(5 downto 0); 
	  rgb : out std_logic_vector(5 downto 0)
	  );
end background_rom;

architecture synth of background_rom is

signal location : std_logic_vector(13 downto 0);
begin
	process (clk) begin
		if rising_edge(clk) then
			case location is
				  when "00000100111100" => rgb <= "100001";
				  when "00000100111101" => rgb <= "100001";
				  when "00000100111110" => rgb <= "100001";
				  when "00000100111111" => rgb <= "100001";
				  when "00000101000000" => rgb <= "100001";
				  when "00000101000001" => rgb <= "100001";
				  when "00000101000010" => rgb <= "100001";
				  when "00000101000101" => rgb <= "100001";
				  when "00000101000110" => rgb <= "100001";
				  when "00000101001010" => rgb <= "100001";
				  when "00000101001011" => rgb <= "100001";
				  when "00000101001110" => rgb <= "100001";
				  when "00000101001111" => rgb <= "100001";
				  when "00000101010000" => rgb <= "100001";
				  when "00000101010001" => rgb <= "100001";
				  when "00000101010101" => rgb <= "100001";
				  when "00000101010110" => rgb <= "100001";
				  when "00000101011000" => rgb <= "100001";
				  when "00000101011001" => rgb <= "100001";
				  when "00000101011010" => rgb <= "100001";
				  when "00000101011110" => rgb <= "100001";
				  when "00000101011111" => rgb <= "100001";
				  when "00000101100000" => rgb <= "100001";
				  when "00000101100001" => rgb <= "100001";
				  when "00001000111100" => rgb <= "100001";
				  when "00001000111101" => rgb <= "100001";
				  when "00001000111110" => rgb <= "100001";
				  when "00001000111111" => rgb <= "100001";
				  when "00001001000000" => rgb <= "100001";
				  when "00001001000001" => rgb <= "100001";
				  when "00001001000010" => rgb <= "100001";
				  when "00001001000101" => rgb <= "100001";
				  when "00001001000110" => rgb <= "100001";
				  when "00001001001010" => rgb <= "100001";
				  when "00001001001011" => rgb <= "100001";
				  when "00001001001110" => rgb <= "100001";
				  when "00001001001111" => rgb <= "100001";
				  when "00001001010000" => rgb <= "100001";
				  when "00001001010001" => rgb <= "100001";
				  when "00001001010101" => rgb <= "100001";
				  when "00001001010110" => rgb <= "100001";
				  when "00001001010111" => rgb <= "100001";
				  when "00001001011000" => rgb <= "100001";
				  when "00001001011001" => rgb <= "100001";
				  when "00001001011110" => rgb <= "100001";
				  when "00001001011111" => rgb <= "100001";
				  when "00001001100000" => rgb <= "100001";
				  when "00001001100001" => rgb <= "100001";
				  when "00001100111111" => rgb <= "100001";
				  when "00001101000000" => rgb <= "100001";
				  when "00001101000101" => rgb <= "100001";
				  when "00001101000110" => rgb <= "100001";
				  when "00001101001010" => rgb <= "100001";
				  when "00001101001011" => rgb <= "100001";
				  when "00001101001110" => rgb <= "100001";
				  when "00001101001111" => rgb <= "100001";
				  when "00001101010101" => rgb <= "100001";
				  when "00001101010110" => rgb <= "100001";
				  when "00001101010111" => rgb <= "100001";
				  when "00001101011000" => rgb <= "100001";
				  when "00001101011110" => rgb <= "100001";
				  when "00001101011111" => rgb <= "100001";
				  when "00010000111111" => rgb <= "100001";
				  when "00010001000000" => rgb <= "100001";
				  when "00010001000101" => rgb <= "100001";
				  when "00010001000110" => rgb <= "100001";
				  when "00010001001010" => rgb <= "100001";
				  when "00010001001011" => rgb <= "100001";
				  when "00010001001110" => rgb <= "100001";
				  when "00010001001111" => rgb <= "100001";
				  when "00010001010000" => rgb <= "100001";
				  when "00010001010001" => rgb <= "100001";
				  when "00010001010101" => rgb <= "100001";
				  when "00010001010110" => rgb <= "100001";
				  when "00010001010111" => rgb <= "100001";
				  when "00010001011000" => rgb <= "100001";
				  when "00010001011110" => rgb <= "100001";
				  when "00010001011111" => rgb <= "100001";
				  when "00010001100000" => rgb <= "100001";
				  when "00010001100001" => rgb <= "100001";
				  when "00010100111111" => rgb <= "100001";
				  when "00010101000000" => rgb <= "100001";
				  when "00010101000101" => rgb <= "100001";
				  when "00010101000110" => rgb <= "100001";
				  when "00010101001010" => rgb <= "100001";
				  when "00010101001011" => rgb <= "100001";
				  when "00010101010000" => rgb <= "100001";
				  when "00010101010001" => rgb <= "100001";
				  when "00010101010101" => rgb <= "100001";
				  when "00010101010110" => rgb <= "100001";
				  when "00010101010111" => rgb <= "100001";
				  when "00010101011000" => rgb <= "100001";
				  when "00010101011001" => rgb <= "100001";
				  when "00010101100000" => rgb <= "100001";
				  when "00010101100001" => rgb <= "100001";
				  when "00011000111111" => rgb <= "100001";
				  when "00011001000000" => rgb <= "100001";
				  when "00011001000101" => rgb <= "100001";
				  when "00011001000110" => rgb <= "100001";
				  when "00011001000111" => rgb <= "100001";
				  when "00011001001000" => rgb <= "100001";
				  when "00011001001001" => rgb <= "100001";
				  when "00011001001010" => rgb <= "100001";
				  when "00011001001011" => rgb <= "100001";
				  when "00011001001110" => rgb <= "100001";
				  when "00011001001111" => rgb <= "100001";
				  when "00011001010000" => rgb <= "100001";
				  when "00011001010001" => rgb <= "100001";
				  when "00011001010101" => rgb <= "100001";
				  when "00011001010110" => rgb <= "100001";
				  when "00011001010111" => rgb <= "100001";
				  when "00011001011000" => rgb <= "100001";
				  when "00011001011001" => rgb <= "100001";
				  when "00011001011010" => rgb <= "100001";
				  when "00011001011110" => rgb <= "100001";
				  when "00011001011111" => rgb <= "100001";
				  when "00011001100000" => rgb <= "100001";
				  when "00011001100001" => rgb <= "100001";
				  when "00011100111111" => rgb <= "100001";
				  when "00011101000000" => rgb <= "100001";
				  when "00011101000110" => rgb <= "100001";
				  when "00011101000111" => rgb <= "100001";
				  when "00011101001000" => rgb <= "100001";
				  when "00011101001001" => rgb <= "100001";
				  when "00011101001010" => rgb <= "100001";
				  when "00011101001110" => rgb <= "100001";
				  when "00011101001111" => rgb <= "100001";
				  when "00011101010000" => rgb <= "100001";
				  when "00011101010001" => rgb <= "100001";
				  when "00011101010101" => rgb <= "100001";
				  when "00011101010110" => rgb <= "100001";
				  when "00011101011000" => rgb <= "100001";
				  when "00011101011001" => rgb <= "100001";
				  when "00011101011010" => rgb <= "100001";
				  when "00011101011110" => rgb <= "100001";
				  when "00011101011111" => rgb <= "100001";
				  when "00011101100000" => rgb <= "100001";
				  when "00011101100001" => rgb <= "100001";
				  when "00101000101001" => rgb <= "111111";
				  when "00101000101010" => rgb <= "111111";
				  when "00101000101011" => rgb <= "111111";
				  when "00101000101101" => rgb <= "111111";
				  when "00101000110000" => rgb <= "111111";
				  when "00101000110001" => rgb <= "111111";
				  when "00101000110010" => rgb <= "111111";
				  when "00101000110100" => rgb <= "111111";
				  when "00101000110110" => rgb <= "111111";
				  when "00101000111000" => rgb <= "111111";
				  when "00101000111001" => rgb <= "111111";
				  when "00101000111011" => rgb <= "111111";
				  when "00101000111100" => rgb <= "111111";
				  when "00101000111101" => rgb <= "111111";
				  when "00101001000000" => rgb <= "111111";
				  when "00101001000001" => rgb <= "111111";
				  when "00101001011101" => rgb <= "111111";
				  when "00101001011110" => rgb <= "111111";
				  when "00101001011111" => rgb <= "111111";
				  when "00101001100001" => rgb <= "111111";
				  when "00101001100100" => rgb <= "111111";
				  when "00101001100101" => rgb <= "111111";
				  when "00101001100110" => rgb <= "111111";
				  when "00101001101000" => rgb <= "111111";
				  when "00101001101010" => rgb <= "111111";
				  when "00101001101100" => rgb <= "111111";
				  when "00101001101101" => rgb <= "111111";
				  when "00101001101111" => rgb <= "111111";
				  when "00101001110000" => rgb <= "111111";
				  when "00101001110001" => rgb <= "111111";
				  when "00101001110100" => rgb <= "111111";
				  when "00101001110101" => rgb <= "111111";
				  when "00101100101001" => rgb <= "111111";
				  when "00101100101011" => rgb <= "111111";
				  when "00101100101101" => rgb <= "111111";
				  when "00101100110000" => rgb <= "111111";
				  when "00101100110010" => rgb <= "111111";
				  when "00101100110100" => rgb <= "111111";
				  when "00101100110110" => rgb <= "111111";
				  when "00101100111000" => rgb <= "111111";
				  when "00101100111011" => rgb <= "111111";
				  when "00101100111101" => rgb <= "111111";
				  when "00101101000001" => rgb <= "111111";
				  when "00101101011101" => rgb <= "111111";
				  when "00101101011111" => rgb <= "111111";
				  when "00101101100001" => rgb <= "111111";
				  when "00101101100100" => rgb <= "111111";
				  when "00101101100110" => rgb <= "111111";
				  when "00101101101000" => rgb <= "111111";
				  when "00101101101010" => rgb <= "111111";
				  when "00101101101100" => rgb <= "111111";
				  when "00101101101111" => rgb <= "111111";
				  when "00101101110001" => rgb <= "111111";
				  when "00101101110011" => rgb <= "111111";
				  when "00101101110110" => rgb <= "111111";
				  when "00110000101001" => rgb <= "111111";
				  when "00110000101010" => rgb <= "111111";
				  when "00110000101011" => rgb <= "111111";
				  when "00110000101101" => rgb <= "111111";
				  when "00110000110000" => rgb <= "111111";
				  when "00110000110001" => rgb <= "111111";
				  when "00110000110010" => rgb <= "111111";
				  when "00110000110101" => rgb <= "111111";
				  when "00110000111000" => rgb <= "111111";
				  when "00110000111001" => rgb <= "111111";
				  when "00110000111011" => rgb <= "111111";
				  when "00110000111100" => rgb <= "111111";
				  when "00110000111101" => rgb <= "111111";
				  when "00110001000001" => rgb <= "111111";
				  when "00110001011101" => rgb <= "111111";
				  when "00110001011110" => rgb <= "111111";
				  when "00110001011111" => rgb <= "111111";
				  when "00110001100001" => rgb <= "111111";
				  when "00110001100100" => rgb <= "111111";
				  when "00110001100101" => rgb <= "111111";
				  when "00110001100110" => rgb <= "111111";
				  when "00110001101001" => rgb <= "111111";
				  when "00110001101100" => rgb <= "111111";
				  when "00110001101101" => rgb <= "111111";
				  when "00110001101111" => rgb <= "111111";
				  when "00110001110000" => rgb <= "111111";
				  when "00110001110001" => rgb <= "111111";
				  when "00110001110101" => rgb <= "111111";
				  when "00110001110110" => rgb <= "111111";
				  when "00110100101001" => rgb <= "111111";
				  when "00110100101101" => rgb <= "111111";
				  when "00110100110000" => rgb <= "111111";
				  when "00110100110010" => rgb <= "111111";
				  when "00110100110101" => rgb <= "111111";
				  when "00110100111000" => rgb <= "111111";
				  when "00110100111011" => rgb <= "111111";
				  when "00110100111100" => rgb <= "111111";
				  when "00110101000001" => rgb <= "111111";
				  when "00110101011101" => rgb <= "111111";
				  when "00110101100001" => rgb <= "111111";
				  when "00110101100100" => rgb <= "111111";
				  when "00110101100110" => rgb <= "111111";
				  when "00110101101001" => rgb <= "111111";
				  when "00110101101100" => rgb <= "111111";
				  when "00110101101111" => rgb <= "111111";
				  when "00110101110000" => rgb <= "111111";
				  when "00110101110100" => rgb <= "111111";
				  when "00111000101001" => rgb <= "111111";
				  when "00111000101101" => rgb <= "111111";
				  when "00111000101110" => rgb <= "111111";
				  when "00111000110000" => rgb <= "111111";
				  when "00111000110010" => rgb <= "111111";
				  when "00111000110101" => rgb <= "111111";
				  when "00111000111000" => rgb <= "111111";
				  when "00111000111001" => rgb <= "111111";
				  when "00111000111011" => rgb <= "111111";
				  when "00111000111101" => rgb <= "111111";
				  when "00111001000000" => rgb <= "111111";
				  when "00111001000001" => rgb <= "111111";
				  when "00111001000010" => rgb <= "111111";
				  when "00111001011101" => rgb <= "111111";
				  when "00111001100001" => rgb <= "111111";
				  when "00111001100010" => rgb <= "111111";
				  when "00111001100100" => rgb <= "111111";
				  when "00111001100110" => rgb <= "111111";
				  when "00111001101001" => rgb <= "111111";
				  when "00111001101100" => rgb <= "111111";
				  when "00111001101101" => rgb <= "111111";
				  when "00111001101111" => rgb <= "111111";
				  when "00111001110001" => rgb <= "111111";
				  when "00111001110100" => rgb <= "111111";
				  when "00111001110101" => rgb <= "111111";
				  when "00111001110110" => rgb <= "111111";
				  when "10000001000000" => rgb <= "111111";
				  when "10000001000001" => rgb <= "111111";
				  when "10000001000010" => rgb <= "111111";
				  when "10000001000011" => rgb <= "111111";
				  when "10000001000100" => rgb <= "111111";
				  when "10000001000101" => rgb <= "111111";
				  when "10000001000110" => rgb <= "111111";
				  when "10000001000111" => rgb <= "111111";
				  when "10000001001000" => rgb <= "111111";
				  when "10000001001001" => rgb <= "111111";
				  when "10000001001010" => rgb <= "111111";
				  when "10000001001011" => rgb <= "111111";
				  when "10000001001100" => rgb <= "111111";
				  when "10000001001101" => rgb <= "111111";
				  when "10000001001110" => rgb <= "111111";
				  when "10000001001111" => rgb <= "111111";
				  when "10000001010000" => rgb <= "111111";
				  when "10000001010001" => rgb <= "111111";
				  when "10000001010010" => rgb <= "111111";
				  when "10000001010011" => rgb <= "111111";
				  when "10000001010100" => rgb <= "111111";
				  when "10000001010101" => rgb <= "111111";
				  when "10000001010110" => rgb <= "111111";
				  when "10000001010111" => rgb <= "111111";
				  when "10000001011000" => rgb <= "111111";
				  when "10000001011001" => rgb <= "111111";
				  when "10000001011010" => rgb <= "111111";
				  when "10000001011011" => rgb <= "111111";
				  when "10000001011100" => rgb <= "111111";
				  when "10000001011101" => rgb <= "111111";
				  when "10000001011110" => rgb <= "111111";
				  when "10000001011111" => rgb <= "111111";
				  when "10000101000000" => rgb <= "111111";
				  when "10000101000001" => rgb <= "111111";
				  when "10000101000010" => rgb <= "111111";
				  when "10000101000011" => rgb <= "111111";
				  when "10000101000100" => rgb <= "111111";
				  when "10000101000101" => rgb <= "111111";
				  when "10000101000110" => rgb <= "111111";
				  when "10000101000111" => rgb <= "111111";
				  when "10000101001000" => rgb <= "111111";
				  when "10000101001001" => rgb <= "111111";
				  when "10000101001010" => rgb <= "111111";
				  when "10000101001011" => rgb <= "111111";
				  when "10000101001100" => rgb <= "111111";
				  when "10000101001101" => rgb <= "111111";
				  when "10000101001110" => rgb <= "111111";
				  when "10000101001111" => rgb <= "111111";
				  when "10000101010000" => rgb <= "111111";
				  when "10000101010001" => rgb <= "111111";
				  when "10000101010010" => rgb <= "111111";
				  when "10000101010011" => rgb <= "111111";
				  when "10000101010100" => rgb <= "111111";
				  when "10000101010101" => rgb <= "111111";
				  when "10000101010110" => rgb <= "111111";
				  when "10000101010111" => rgb <= "111111";
				  when "10000101011000" => rgb <= "111111";
				  when "10000101011001" => rgb <= "111111";
				  when "10000101011010" => rgb <= "111111";
				  when "10000101011011" => rgb <= "111111";
				  when "10000101011100" => rgb <= "111111";
				  when "10000101011101" => rgb <= "111111";
				  when "10000101011110" => rgb <= "111111";
				  when "10000101011111" => rgb <= "111111";
				  when "10001001000000" => rgb <= "111111";
				  when "10001001000001" => rgb <= "111111";
				  when "10001001000010" => rgb <= "111111";
				  when "10001001000011" => rgb <= "111111";
				  when "10001001000100" => rgb <= "111111";
				  when "10001001000101" => rgb <= "111111";
				  when "10001001000110" => rgb <= "111111";
				  when "10001001000111" => rgb <= "111111";
				  when "10001001001000" => rgb <= "111111";
				  when "10001001001001" => rgb <= "111111";
				  when "10001001001010" => rgb <= "111111";
				  when "10001001001011" => rgb <= "111111";
				  when "10001001001100" => rgb <= "111111";
				  when "10001001001101" => rgb <= "111111";
				  when "10001001001110" => rgb <= "111111";
				  when "10001001001111" => rgb <= "111111";
				  when "10001001010000" => rgb <= "111111";
				  when "10001001010001" => rgb <= "111111";
				  when "10001001010010" => rgb <= "111111";
				  when "10001001010011" => rgb <= "111111";
				  when "10001001010100" => rgb <= "111111";
				  when "10001001010101" => rgb <= "111111";
				  when "10001001010110" => rgb <= "111111";
				  when "10001001010111" => rgb <= "111111";
				  when "10001001011000" => rgb <= "111111";
				  when "10001001011001" => rgb <= "111111";
				  when "10001001011010" => rgb <= "111111";
				  when "10001001011011" => rgb <= "111111";
				  when "10001001011100" => rgb <= "111111";
				  when "10001001011101" => rgb <= "111111";
				  when "10001001011110" => rgb <= "111111";
				  when "10001001011111" => rgb <= "111111";
				  when "10001101000000" => rgb <= "111111";
				  when "10001101000001" => rgb <= "111111";
				  when "10001101000010" => rgb <= "111111";
				  when "10001101000011" => rgb <= "111111";
				  when "10001101000100" => rgb <= "111111";
				  when "10001101000101" => rgb <= "111111";
				  when "10001101000110" => rgb <= "111111";
				  when "10001101000111" => rgb <= "111111";
				  when "10001101001000" => rgb <= "111111";
				  when "10001101001001" => rgb <= "111111";
				  when "10001101001010" => rgb <= "111111";
				  when "10001101001011" => rgb <= "111111";
				  when "10001101001100" => rgb <= "111111";
				  when "10001101001101" => rgb <= "111111";
				  when "10001101001110" => rgb <= "111111";
				  when "10001101001111" => rgb <= "111111";
				  when "10001101010000" => rgb <= "111111";
				  when "10001101010001" => rgb <= "111111";
				  when "10001101010010" => rgb <= "111111";
				  when "10001101010011" => rgb <= "111111";
				  when "10001101010100" => rgb <= "111111";
				  when "10001101010101" => rgb <= "111111";
				  when "10001101010110" => rgb <= "111111";
				  when "10001101010111" => rgb <= "111111";
				  when "10001101011000" => rgb <= "111111";
				  when "10001101011001" => rgb <= "111111";
				  when "10001101011010" => rgb <= "111111";
				  when "10001101011011" => rgb <= "111111";
				  when "10001101011100" => rgb <= "111111";
				  when "10001101011101" => rgb <= "111111";
				  when "10001101011110" => rgb <= "111111";
				  when "10001101011111" => rgb <= "111111";
				  when "10010001000000" => rgb <= "111111";
				  when "10010001000001" => rgb <= "111111";
				  when "10010001000100" => rgb <= "111111";
				  when "10010001000101" => rgb <= "111111";
				  when "10010001001000" => rgb <= "111111";
				  when "10010001001001" => rgb <= "111111";
				  when "10010001001100" => rgb <= "111111";
				  when "10010001001101" => rgb <= "111111";
				  when "10010001001110" => rgb <= "111111";
				  when "10010001010001" => rgb <= "111111";
				  when "10010001010010" => rgb <= "111111";
				  when "10010001010011" => rgb <= "111111";
				  when "10010001010110" => rgb <= "111111";
				  when "10010001010111" => rgb <= "111111";
				  when "10010001011010" => rgb <= "111111";
				  when "10010001011011" => rgb <= "111111";
				  when "10010001011110" => rgb <= "111111";
				  when "10010001011111" => rgb <= "111111";
				  when "10010101000000" => rgb <= "111111";
				  when "10010101000001" => rgb <= "111111";
				  when "10010101000100" => rgb <= "111111";
				  when "10010101000101" => rgb <= "111111";
				  when "10010101001000" => rgb <= "111111";
				  when "10010101001001" => rgb <= "111111";
				  when "10010101001100" => rgb <= "111111";
				  when "10010101001101" => rgb <= "111111";
				  when "10010101001110" => rgb <= "111111";
				  when "10010101010001" => rgb <= "111111";
				  when "10010101010010" => rgb <= "111111";
				  when "10010101010011" => rgb <= "111111";
				  when "10010101010110" => rgb <= "111111";
				  when "10010101010111" => rgb <= "111111";
				  when "10010101011010" => rgb <= "111111";
				  when "10010101011011" => rgb <= "111111";
				  when "10010101011110" => rgb <= "111111";
				  when "10010101011111" => rgb <= "111111";
				  when "10011001000000" => rgb <= "111111";
				  when "10011001000001" => rgb <= "111111";
				  when "10011001000100" => rgb <= "111111";
				  when "10011001000101" => rgb <= "111111";
				  when "10011001001000" => rgb <= "111111";
				  when "10011001001001" => rgb <= "111111";
				  when "10011001001100" => rgb <= "111111";
				  when "10011001001101" => rgb <= "111111";
				  when "10011001001110" => rgb <= "111111";
				  when "10011001010001" => rgb <= "111111";
				  when "10011001010010" => rgb <= "111111";
				  when "10011001010011" => rgb <= "111111";
				  when "10011001010110" => rgb <= "111111";
				  when "10011001010111" => rgb <= "111111";
				  when "10011001011010" => rgb <= "111111";
				  when "10011001011011" => rgb <= "111111";
				  when "10011001011110" => rgb <= "111111";
				  when "10011001011111" => rgb <= "111111";
				  when "10011101000000" => rgb <= "111111";
				  when "10011101000001" => rgb <= "111111";
				  when "10011101000100" => rgb <= "111111";
				  when "10011101000101" => rgb <= "111111";
				  when "10011101001000" => rgb <= "111111";
				  when "10011101001001" => rgb <= "111111";
				  when "10011101001100" => rgb <= "111111";
				  when "10011101001101" => rgb <= "111111";
				  when "10011101001110" => rgb <= "111111";
				  when "10011101010001" => rgb <= "111111";
				  when "10011101010010" => rgb <= "111111";
				  when "10011101010011" => rgb <= "111111";
				  when "10011101010110" => rgb <= "111111";
				  when "10011101010111" => rgb <= "111111";
				  when "10011101011010" => rgb <= "111111";
				  when "10011101011011" => rgb <= "111111";
				  when "10011101011110" => rgb <= "111111";
				  when "10011101011111" => rgb <= "111111";
				  when "10100001000000" => rgb <= "111111";
				  when "10100001000001" => rgb <= "111111";
				  when "10100001000100" => rgb <= "111111";
				  when "10100001000101" => rgb <= "111111";
				  when "10100001001000" => rgb <= "111111";
				  when "10100001001001" => rgb <= "111111";
				  when "10100001001100" => rgb <= "111111";
				  when "10100001001101" => rgb <= "111111";
				  when "10100001001110" => rgb <= "111111";
				  when "10100001010001" => rgb <= "111111";
				  when "10100001010010" => rgb <= "111111";
				  when "10100001010011" => rgb <= "111111";
				  when "10100001010110" => rgb <= "111111";
				  when "10100001010111" => rgb <= "111111";
				  when "10100001011010" => rgb <= "111111";
				  when "10100001011011" => rgb <= "111111";
				  when "10100001011110" => rgb <= "111111";
				  when "10100001011111" => rgb <= "111111";
				  when "10100101000000" => rgb <= "111111";
				  when "10100101000001" => rgb <= "111111";
				  when "10100101000100" => rgb <= "111111";
				  when "10100101000101" => rgb <= "111111";
				  when "10100101001000" => rgb <= "111111";
				  when "10100101001001" => rgb <= "111111";
				  when "10100101001100" => rgb <= "111111";
				  when "10100101001101" => rgb <= "111111";
				  when "10100101001110" => rgb <= "111111";
				  when "10100101010001" => rgb <= "111111";
				  when "10100101010010" => rgb <= "111111";
				  when "10100101010011" => rgb <= "111111";
				  when "10100101010110" => rgb <= "111111";
				  when "10100101010111" => rgb <= "111111";
				  when "10100101011010" => rgb <= "111111";
				  when "10100101011011" => rgb <= "111111";
				  when "10100101011110" => rgb <= "111111";
				  when "10100101011111" => rgb <= "111111";
				  when "10101001000000" => rgb <= "111111";
				  when "10101001000001" => rgb <= "111111";
				  when "10101001000010" => rgb <= "111111";
				  when "10101001000011" => rgb <= "111111";
				  when "10101001000100" => rgb <= "111111";
				  when "10101001000101" => rgb <= "111111";
				  when "10101001000110" => rgb <= "111111";
				  when "10101001000111" => rgb <= "111111";
				  when "10101001001000" => rgb <= "111111";
				  when "10101001001001" => rgb <= "111111";
				  when "10101001001010" => rgb <= "111111";
				  when "10101001001011" => rgb <= "111111";
				  when "10101001001100" => rgb <= "111111";
				  when "10101001001101" => rgb <= "111111";
				  when "10101001001110" => rgb <= "111111";
				  when "10101001001111" => rgb <= "111111";
				  when "10101001010000" => rgb <= "111111";
				  when "10101001010001" => rgb <= "111111";
				  when "10101001010010" => rgb <= "111111";
				  when "10101001010011" => rgb <= "111111";
				  when "10101001010100" => rgb <= "111111";
				  when "10101001010101" => rgb <= "111111";
				  when "10101001010110" => rgb <= "111111";
				  when "10101001010111" => rgb <= "111111";
				  when "10101001011000" => rgb <= "111111";
				  when "10101001011001" => rgb <= "111111";
				  when "10101001011010" => rgb <= "111111";
				  when "10101001011011" => rgb <= "111111";
				  when "10101001011100" => rgb <= "111111";
				  when "10101001011101" => rgb <= "111111";
				  when "10101001011110" => rgb <= "111111";
				  when "10101001011111" => rgb <= "111111";
				  when "10101101000000" => rgb <= "111111";
				  when "10101101000001" => rgb <= "111111";
				  when "10101101000010" => rgb <= "111111";
				  when "10101101000011" => rgb <= "111111";
				  when "10101101000100" => rgb <= "111111";
				  when "10101101000101" => rgb <= "111111";
				  when "10101101000110" => rgb <= "111111";
				  when "10101101000111" => rgb <= "111111";
				  when "10101101001000" => rgb <= "111111";
				  when "10101101001001" => rgb <= "111111";
				  when "10101101001010" => rgb <= "111111";
				  when "10101101001011" => rgb <= "111111";
				  when "10101101001100" => rgb <= "111111";
				  when "10101101001101" => rgb <= "111111";
				  when "10101101001110" => rgb <= "111111";
				  when "10101101001111" => rgb <= "111111";
				  when "10101101010000" => rgb <= "111111";
				  when "10101101010001" => rgb <= "111111";
				  when "10101101010010" => rgb <= "111111";
				  when "10101101010011" => rgb <= "111111";
				  when "10101101010100" => rgb <= "111111";
				  when "10101101010101" => rgb <= "111111";
				  when "10101101010110" => rgb <= "111111";
				  when "10101101010111" => rgb <= "111111";
				  when "10101101011000" => rgb <= "111111";
				  when "10101101011001" => rgb <= "111111";
				  when "10101101011010" => rgb <= "111111";
				  when "10101101011011" => rgb <= "111111";
				  when "10101101011100" => rgb <= "111111";
				  when "10101101011101" => rgb <= "111111";
				  when "10101101011110" => rgb <= "111111";
				  when "10101101011111" => rgb <= "111111";
				  when "10110001000000" => rgb <= "111111";
				  when "10110001000001" => rgb <= "111111";
				  when "10110001000010" => rgb <= "111111";
				  when "10110001000011" => rgb <= "111111";
				  when "10110001000100" => rgb <= "111111";
				  when "10110001000101" => rgb <= "111111";
				  when "10110001000110" => rgb <= "111111";
				  when "10110001000111" => rgb <= "111111";
				  when "10110001001000" => rgb <= "111111";
				  when "10110001001001" => rgb <= "111111";
				  when "10110001001010" => rgb <= "111111";
				  when "10110001001011" => rgb <= "111111";
				  when "10110001001100" => rgb <= "111111";
				  when "10110001001101" => rgb <= "111111";
				  when "10110001001110" => rgb <= "111111";
				  when "10110001001111" => rgb <= "111111";
				  when "10110001010000" => rgb <= "111111";
				  when "10110001010001" => rgb <= "111111";
				  when "10110001010010" => rgb <= "111111";
				  when "10110001010011" => rgb <= "111111";
				  when "10110001010100" => rgb <= "111111";
				  when "10110001010101" => rgb <= "111111";
				  when "10110001010110" => rgb <= "111111";
				  when "10110001010111" => rgb <= "111111";
				  when "10110001011000" => rgb <= "111111";
				  when "10110001011001" => rgb <= "111111";
				  when "10110001011010" => rgb <= "111111";
				  when "10110001011011" => rgb <= "111111";
				  when "10110001011100" => rgb <= "111111";
				  when "10110001011101" => rgb <= "111111";
				  when "10110001011110" => rgb <= "111111";
				  when "10110001011111" => rgb <= "111111";
				  when "10110101000000" => rgb <= "111111";
				  when "10110101000001" => rgb <= "111111";
				  when "10110101000010" => rgb <= "111111";
				  when "10110101000011" => rgb <= "111111";
				  when "10110101000100" => rgb <= "111111";
				  when "10110101000101" => rgb <= "111111";
				  when "10110101000110" => rgb <= "111111";
				  when "10110101000111" => rgb <= "111111";
				  when "10110101001000" => rgb <= "111111";
				  when "10110101001001" => rgb <= "111111";
				  when "10110101001010" => rgb <= "111111";
				  when "10110101001011" => rgb <= "111111";
				  when "10110101001100" => rgb <= "111111";
				  when "10110101001101" => rgb <= "111111";
				  when "10110101001110" => rgb <= "111111";
				  when "10110101001111" => rgb <= "111111";
				  when "10110101010000" => rgb <= "111111";
				  when "10110101010001" => rgb <= "111111";
				  when "10110101010010" => rgb <= "111111";
				  when "10110101010011" => rgb <= "111111";
				  when "10110101010100" => rgb <= "111111";
				  when "10110101010101" => rgb <= "111111";
				  when "10110101010110" => rgb <= "111111";
				  when "10110101010111" => rgb <= "111111";
				  when "10110101011000" => rgb <= "111111";
				  when "10110101011001" => rgb <= "111111";
				  when "10110101011010" => rgb <= "111111";
				  when "10110101011011" => rgb <= "111111";
				  when "10110101011100" => rgb <= "111111";
				  when "10110101011101" => rgb <= "111111";
				  when "10110101011110" => rgb <= "111111";
				  when "10110101011111" => rgb <= "111111";
				  when "10111001000000" => rgb <= "111111";
				  when "10111001000001" => rgb <= "111111";
				  when "10111001000110" => rgb <= "111111";
				  when "10111001000111" => rgb <= "111111";
				  when "10111001001000" => rgb <= "111111";
				  when "10111001001001" => rgb <= "111111";
				  when "10111001001010" => rgb <= "111111";
				  when "10111001001011" => rgb <= "111111";
				  when "10111001001100" => rgb <= "111111";
				  when "10111001001101" => rgb <= "111111";
				  when "10111001010010" => rgb <= "111111";
				  when "10111001010011" => rgb <= "111111";
				  when "10111001011000" => rgb <= "111111";
				  when "10111001011001" => rgb <= "111111";
				  when "10111001011110" => rgb <= "111111";
				  when "10111001011111" => rgb <= "111111";
				  when "10111101000000" => rgb <= "111111";
				  when "10111101000001" => rgb <= "111111";
				  when "10111101000110" => rgb <= "111111";
				  when "10111101000111" => rgb <= "111111";
				  when "10111101001000" => rgb <= "111111";
				  when "10111101001001" => rgb <= "111111";
				  when "10111101001010" => rgb <= "111111";
				  when "10111101001011" => rgb <= "111111";
				  when "10111101001100" => rgb <= "111111";
				  when "10111101001101" => rgb <= "111111";
				  when "10111101010010" => rgb <= "111111";
				  when "10111101010011" => rgb <= "111111";
				  when "10111101011000" => rgb <= "111111";
				  when "10111101011001" => rgb <= "111111";
				  when "10111101011110" => rgb <= "111111";
				  when "10111101011111" => rgb <= "111111";
				  when "11000001000000" => rgb <= "111111";
				  when "11000001000001" => rgb <= "111111";
				  when "11000001000110" => rgb <= "111111";
				  when "11000001000111" => rgb <= "111111";
				  when "11000001001000" => rgb <= "111111";
				  when "11000001001001" => rgb <= "111111";
				  when "11000001001010" => rgb <= "001011";
				  when "11000001001011" => rgb <= "001011";
				  when "11000001001100" => rgb <= "111111";
				  when "11000001001101" => rgb <= "111111";
				  when "11000001001110" => rgb <= "111111";
				  when "11000001001111" => rgb <= "111111";
				  when "11000001010000" => rgb <= "111111";
				  when "11000001010001" => rgb <= "111111";
				  when "11000001010010" => rgb <= "111111";
				  when "11000001010011" => rgb <= "111111";
				  when "11000001010100" => rgb <= "111111";
				  when "11000001010101" => rgb <= "111111";
				  when "11000001010110" => rgb <= "111111";
				  when "11000001010111" => rgb <= "111111";
				  when "11000001011000" => rgb <= "111111";
				  when "11000001011001" => rgb <= "111111";
				  when "11000001011010" => rgb <= "111111";
				  when "11000001011011" => rgb <= "111111";
				  when "11000001011100" => rgb <= "111111";
				  when "11000001011101" => rgb <= "111111";
				  when "11000001011110" => rgb <= "111111";
				  when "11000001011111" => rgb <= "111111";
				  when "11000101000000" => rgb <= "111111";
				  when "11000101000001" => rgb <= "111111";
				  when "11000101000110" => rgb <= "111111";
				  when "11000101000111" => rgb <= "111111";
				  when "11000101001000" => rgb <= "111111";
				  when "11000101001001" => rgb <= "111111";
				  when "11000101001010" => rgb <= "001011";
				  when "11000101001011" => rgb <= "001011";
				  when "11000101001100" => rgb <= "111111";
				  when "11000101001101" => rgb <= "111111";
				  when "11000101001110" => rgb <= "111111";
				  when "11000101001111" => rgb <= "111111";
				  when "11000101010000" => rgb <= "111111";
				  when "11000101010001" => rgb <= "111111";
				  when "11000101010010" => rgb <= "111111";
				  when "11000101010011" => rgb <= "111111";
				  when "11000101010100" => rgb <= "111111";
				  when "11000101010101" => rgb <= "111111";
				  when "11000101010110" => rgb <= "111111";
				  when "11000101010111" => rgb <= "111111";
				  when "11000101011000" => rgb <= "111111";
				  when "11000101011001" => rgb <= "111111";
				  when "11000101011010" => rgb <= "111111";
				  when "11000101011011" => rgb <= "111111";
				  when "11000101011100" => rgb <= "111111";
				  when "11000101011101" => rgb <= "111111";
				  when "11000101011110" => rgb <= "111111";
				  when "11000101011111" => rgb <= "111111";
				  when "11001001000000" => rgb <= "111111";
				  when "11001001000001" => rgb <= "111111";
				  when "11001001000010" => rgb <= "111111";
				  when "11001001000011" => rgb <= "111111";
				  when "11001001000100" => rgb <= "111111";
				  when "11001001000101" => rgb <= "111111";
				  when "11001001000110" => rgb <= "111111";
				  when "11001001000111" => rgb <= "111111";
				  when "11001001001000" => rgb <= "111111";
				  when "11001001001001" => rgb <= "111111";
				  when "11001001001010" => rgb <= "001011";
				  when "11001001001011" => rgb <= "001011";
				  when "11001001001100" => rgb <= "111111";
				  when "11001001001101" => rgb <= "111111";
				  when "11001001001110" => rgb <= "111111";
				  when "11001001001111" => rgb <= "111111";
				  when "11001001010000" => rgb <= "111111";
				  when "11001001010001" => rgb <= "111111";
				  when "11001001010010" => rgb <= "111111";
				  when "11001001010011" => rgb <= "111111";
				  when "11001001010100" => rgb <= "111111";
				  when "11001001010101" => rgb <= "111111";
				  when "11001001010110" => rgb <= "111111";
				  when "11001001010111" => rgb <= "111111";
				  when "11001001011000" => rgb <= "111111";
				  when "11001001011001" => rgb <= "111111";
				  when "11001001011010" => rgb <= "111111";
				  when "11001001011011" => rgb <= "111111";
				  when "11001001011100" => rgb <= "111111";
				  when "11001001011101" => rgb <= "111111";
				  when "11001001011110" => rgb <= "111111";
				  when "11001001011111" => rgb <= "111111";
				  when "11001101000000" => rgb <= "111111";
				  when "11001101000001" => rgb <= "111111";
				  when "11001101000010" => rgb <= "111111";
				  when "11001101000011" => rgb <= "111111";
				  when "11001101000100" => rgb <= "111111";
				  when "11001101000101" => rgb <= "111111";
				  when "11001101000110" => rgb <= "111111";
				  when "11001101000111" => rgb <= "111111";
				  when "11001101001000" => rgb <= "111111";
				  when "11001101001001" => rgb <= "111111";
				  when "11001101001010" => rgb <= "001011";
				  when "11001101001011" => rgb <= "001011";
				  when "11001101001100" => rgb <= "111111";
				  when "11001101001101" => rgb <= "111111";
				  when "11001101001110" => rgb <= "111111";
				  when "11001101001111" => rgb <= "111111";
				  when "11001101010000" => rgb <= "111111";
				  when "11001101010001" => rgb <= "111111";
				  when "11001101010010" => rgb <= "111111";
				  when "11001101010011" => rgb <= "111111";
				  when "11001101010100" => rgb <= "111111";
				  when "11001101010101" => rgb <= "111111";
				  when "11001101010110" => rgb <= "111111";
				  when "11001101010111" => rgb <= "111111";
				  when "11001101011000" => rgb <= "111111";
				  when "11001101011001" => rgb <= "111111";
				  when "11001101011010" => rgb <= "111111";
				  when "11001101011011" => rgb <= "111111";
				  when "11001101011100" => rgb <= "111111";
				  when "11001101011101" => rgb <= "111111";
				  when "11001101011110" => rgb <= "111111";
				  when "11001101011111" => rgb <= "111111";
				  when "11010000000000" => rgb <= "111111";
				  when "11010000000001" => rgb <= "111111";
				  when "11010000000010" => rgb <= "111111";
				  when "11010000000011" => rgb <= "111111";
				  when "11010000000100" => rgb <= "111111";
				  when "11010000000101" => rgb <= "111111";
				  when "11010000000110" => rgb <= "111111";
				  when "11010000000111" => rgb <= "111111";
				  when "11010000001000" => rgb <= "111111";
				  when "11010000001001" => rgb <= "111111";
				  when "11010000001010" => rgb <= "111111";
				  when "11010000001011" => rgb <= "111111";
				  when "11010000001100" => rgb <= "111111";
				  when "11010000001101" => rgb <= "111111";
				  when "11010000001110" => rgb <= "111111";
				  when "11010000001111" => rgb <= "111111";
				  when "11010000010000" => rgb <= "111111";
				  when "11010000010001" => rgb <= "111111";
				  when "11010000010010" => rgb <= "111111";
				  when "11010000010011" => rgb <= "111111";
				  when "11010000010100" => rgb <= "111111";
				  when "11010000010101" => rgb <= "111111";
				  when "11010000010110" => rgb <= "111111";
				  when "11010000010111" => rgb <= "111111";
				  when "11010000011000" => rgb <= "111111";
				  when "11010000011001" => rgb <= "111111";
				  when "11010000011010" => rgb <= "111111";
				  when "11010000011011" => rgb <= "111111";
				  when "11010000011100" => rgb <= "111111";
				  when "11010000011101" => rgb <= "111111";
				  when "11010000011110" => rgb <= "111111";
				  when "11010000011111" => rgb <= "111111";
				  when "11010000100000" => rgb <= "111111";
				  when "11010000100001" => rgb <= "111111";
				  when "11010000100010" => rgb <= "111111";
				  when "11010000100011" => rgb <= "111111";
				  when "11010000100100" => rgb <= "111111";
				  when "11010000100101" => rgb <= "111111";
				  when "11010000100110" => rgb <= "111111";
				  when "11010000100111" => rgb <= "111111";
				  when "11010000101000" => rgb <= "111111";
				  when "11010000101001" => rgb <= "111111";
				  when "11010000101010" => rgb <= "111111";
				  when "11010000101011" => rgb <= "111111";
				  when "11010000101100" => rgb <= "111111";
				  when "11010000101101" => rgb <= "111111";
				  when "11010000101110" => rgb <= "111111";
				  when "11010000101111" => rgb <= "111111";
				  when "11010000110000" => rgb <= "111111";
				  when "11010000110001" => rgb <= "111111";
				  when "11010000110010" => rgb <= "111111";
				  when "11010000110011" => rgb <= "111111";
				  when "11010000110100" => rgb <= "111111";
				  when "11010000110101" => rgb <= "111111";
				  when "11010000110110" => rgb <= "111111";
				  when "11010000110111" => rgb <= "111111";
				  when "11010000111000" => rgb <= "111111";
				  when "11010000111001" => rgb <= "111111";
				  when "11010000111010" => rgb <= "111111";
				  when "11010000111011" => rgb <= "111111";
				  when "11010000111100" => rgb <= "111111";
				  when "11010000111101" => rgb <= "111111";
				  when "11010000111110" => rgb <= "111111";
				  when "11010000111111" => rgb <= "111111";
				  when "11010001000000" => rgb <= "111111";
				  when "11010001000001" => rgb <= "111111";
				  when "11010001000010" => rgb <= "111111";
				  when "11010001000011" => rgb <= "111111";
				  when "11010001000100" => rgb <= "111111";
				  when "11010001000101" => rgb <= "111111";
				  when "11010001000110" => rgb <= "111111";
				  when "11010001000111" => rgb <= "111111";
				  when "11010001001000" => rgb <= "111111";
				  when "11010001001001" => rgb <= "111111";
				  when "11010001001010" => rgb <= "111111";
				  when "11010001001011" => rgb <= "111111";
				  when "11010001001100" => rgb <= "111111";
				  when "11010001001101" => rgb <= "111111";
				  when "11010001001110" => rgb <= "111111";
				  when "11010001001111" => rgb <= "111111";
				  when "11010001010000" => rgb <= "111111";
				  when "11010001010001" => rgb <= "111111";
				  when "11010001010010" => rgb <= "111111";
				  when "11010001010011" => rgb <= "111111";
				  when "11010001010100" => rgb <= "111111";
				  when "11010001010101" => rgb <= "111111";
				  when "11010001010110" => rgb <= "111111";
				  when "11010001010111" => rgb <= "111111";
				  when "11010001011000" => rgb <= "111111";
				  when "11010001011001" => rgb <= "111111";
				  when "11010001011010" => rgb <= "111111";
				  when "11010001011011" => rgb <= "111111";
				  when "11010001011100" => rgb <= "111111";
				  when "11010001011101" => rgb <= "111111";
				  when "11010001011110" => rgb <= "111111";
				  when "11010001011111" => rgb <= "111111";
				  when "11010001100000" => rgb <= "111111";
				  when "11010001100001" => rgb <= "111111";
				  when "11010001100010" => rgb <= "111111";
				  when "11010001100011" => rgb <= "111111";
				  when "11010001100100" => rgb <= "111111";
				  when "11010001100101" => rgb <= "111111";
				  when "11010001100110" => rgb <= "111111";
				  when "11010001100111" => rgb <= "111111";
				  when "11010001101000" => rgb <= "111111";
				  when "11010001101001" => rgb <= "111111";
				  when "11010001101010" => rgb <= "111111";
				  when "11010001101011" => rgb <= "111111";
				  when "11010001101100" => rgb <= "111111";
				  when "11010001101101" => rgb <= "111111";
				  when "11010001101110" => rgb <= "111111";
				  when "11010001101111" => rgb <= "111111";
				  when "11010001110000" => rgb <= "111111";
				  when "11010001110001" => rgb <= "111111";
				  when "11010001110010" => rgb <= "111111";
				  when "11010001110011" => rgb <= "111111";
				  when "11010001110100" => rgb <= "111111";
				  when "11010001110101" => rgb <= "111111";
				  when "11010001110110" => rgb <= "111111";
				  when "11010001110111" => rgb <= "111111";
				  when "11010001111000" => rgb <= "111111";
				  when "11010001111001" => rgb <= "111111";
				  when "11010001111010" => rgb <= "111111";
				  when "11010001111011" => rgb <= "111111";
				  when "11010001111100" => rgb <= "111111";
				  when "11010001111101" => rgb <= "111111";
				  when "11010001111110" => rgb <= "111111";
				  when "11010001111111" => rgb <= "111111";
				  when "11010010000000" => rgb <= "111111";
				  when "11010010000001" => rgb <= "111111";
				  when "11010010000010" => rgb <= "111111";
				  when "11010010000011" => rgb <= "111111";
				  when "11010010000100" => rgb <= "111111";
				  when "11010010000101" => rgb <= "111111";
				  when "11010010000110" => rgb <= "111111";
				  when "11010010000111" => rgb <= "111111";
				  when "11010010001000" => rgb <= "111111";
				  when "11010010001001" => rgb <= "111111";
				  when "11010010001010" => rgb <= "111111";
				  when "11010010001011" => rgb <= "111111";
				  when "11010010001100" => rgb <= "111111";
				  when "11010010001101" => rgb <= "111111";
				  when "11010010001110" => rgb <= "111111";
				  when "11010010001111" => rgb <= "111111";
				  when "11010010010000" => rgb <= "111111";
				  when "11010010010001" => rgb <= "111111";
				  when "11010010010010" => rgb <= "111111";
				  when "11010010010011" => rgb <= "111111";
				  when "11010010010100" => rgb <= "111111";
				  when "11010010010101" => rgb <= "111111";
				  when "11010010010110" => rgb <= "111111";
				  when "11010010010111" => rgb <= "111111";
				  when "11010010011000" => rgb <= "111111";
				  when "11010010011001" => rgb <= "111111";
				  when "11010010011010" => rgb <= "111111";
				  when "11010010011011" => rgb <= "111111";
				  when "11010010011100" => rgb <= "111111";
				  when "11010010011101" => rgb <= "111111";
				  when "11010010011110" => rgb <= "111111";
				  when "11010010011111" => rgb <= "111111";
				  when "11010100000000" => rgb <= "111111";
				  when "11010100000001" => rgb <= "111111";
				  when "11010100000010" => rgb <= "111111";
				  when "11010100000011" => rgb <= "111111";
				  when "11010100000100" => rgb <= "111111";
				  when "11010100000101" => rgb <= "111111";
				  when "11010100000110" => rgb <= "111111";
				  when "11010100000111" => rgb <= "111111";
				  when "11010100001000" => rgb <= "111111";
				  when "11010100001001" => rgb <= "111111";
				  when "11010100001010" => rgb <= "111111";
				  when "11010100001011" => rgb <= "111111";
				  when "11010100001100" => rgb <= "111111";
				  when "11010100001101" => rgb <= "111111";
				  when "11010100001110" => rgb <= "111111";
				  when "11010100001111" => rgb <= "111111";
				  when "11010100010000" => rgb <= "111111";
				  when "11010100010001" => rgb <= "111111";
				  when "11010100010010" => rgb <= "111111";
				  when "11010100010011" => rgb <= "111111";
				  when "11010100010100" => rgb <= "111111";
				  when "11010100010101" => rgb <= "111111";
				  when "11010100010110" => rgb <= "111111";
				  when "11010100010111" => rgb <= "111111";
				  when "11010100011000" => rgb <= "111111";
				  when "11010100011001" => rgb <= "111111";
				  when "11010100011010" => rgb <= "111111";
				  when "11010100011011" => rgb <= "111111";
				  when "11010100011100" => rgb <= "111111";
				  when "11010100011101" => rgb <= "111111";
				  when "11010100011110" => rgb <= "111111";
				  when "11010100011111" => rgb <= "111111";
				  when "11010100100000" => rgb <= "111111";
				  when "11010100100001" => rgb <= "111111";
				  when "11010100100010" => rgb <= "111111";
				  when "11010100100011" => rgb <= "111111";
				  when "11010100100100" => rgb <= "111111";
				  when "11010100100101" => rgb <= "111111";
				  when "11010100100110" => rgb <= "111111";
				  when "11010100100111" => rgb <= "111111";
				  when "11010100101000" => rgb <= "111111";
				  when "11010100101001" => rgb <= "111111";
				  when "11010100101010" => rgb <= "111111";
				  when "11010100101011" => rgb <= "111111";
				  when "11010100101100" => rgb <= "111111";
				  when "11010100101101" => rgb <= "111111";
				  when "11010100101110" => rgb <= "111111";
				  when "11010100101111" => rgb <= "111111";
				  when "11010100110000" => rgb <= "111111";
				  when "11010100110001" => rgb <= "111111";
				  when "11010100110010" => rgb <= "111111";
				  when "11010100110011" => rgb <= "111111";
				  when "11010100110100" => rgb <= "111111";
				  when "11010100110101" => rgb <= "111111";
				  when "11010100110110" => rgb <= "111111";
				  when "11010100110111" => rgb <= "111111";
				  when "11010100111000" => rgb <= "111111";
				  when "11010100111001" => rgb <= "111111";
				  when "11010100111010" => rgb <= "111111";
				  when "11010100111011" => rgb <= "111111";
				  when "11010100111100" => rgb <= "111111";
				  when "11010100111101" => rgb <= "111111";
				  when "11010100111110" => rgb <= "111111";
				  when "11010100111111" => rgb <= "111111";
				  when "11010101000000" => rgb <= "111111";
				  when "11010101000001" => rgb <= "111111";
				  when "11010101000010" => rgb <= "111111";
				  when "11010101000011" => rgb <= "111111";
				  when "11010101000100" => rgb <= "111111";
				  when "11010101000101" => rgb <= "111111";
				  when "11010101000110" => rgb <= "111111";
				  when "11010101000111" => rgb <= "111111";
				  when "11010101001000" => rgb <= "111111";
				  when "11010101001001" => rgb <= "111111";
				  when "11010101001010" => rgb <= "111111";
				  when "11010101001011" => rgb <= "111111";
				  when "11010101001100" => rgb <= "111111";
				  when "11010101001101" => rgb <= "111111";
				  when "11010101001110" => rgb <= "111111";
				  when "11010101001111" => rgb <= "111111";
				  when "11010101010000" => rgb <= "111111";
				  when "11010101010001" => rgb <= "111111";
				  when "11010101010010" => rgb <= "111111";
				  when "11010101010011" => rgb <= "111111";
				  when "11010101010100" => rgb <= "111111";
				  when "11010101010101" => rgb <= "111111";
				  when "11010101010110" => rgb <= "111111";
				  when "11010101010111" => rgb <= "111111";
				  when "11010101011000" => rgb <= "111111";
				  when "11010101011001" => rgb <= "111111";
				  when "11010101011010" => rgb <= "111111";
				  when "11010101011011" => rgb <= "111111";
				  when "11010101011100" => rgb <= "111111";
				  when "11010101011101" => rgb <= "111111";
				  when "11010101011110" => rgb <= "111111";
				  when "11010101011111" => rgb <= "111111";
				  when "11010101100000" => rgb <= "111111";
				  when "11010101100001" => rgb <= "111111";
				  when "11010101100010" => rgb <= "111111";
				  when "11010101100011" => rgb <= "111111";
				  when "11010101100100" => rgb <= "111111";
				  when "11010101100101" => rgb <= "111111";
				  when "11010101100110" => rgb <= "111111";
				  when "11010101100111" => rgb <= "111111";
				  when "11010101101000" => rgb <= "111111";
				  when "11010101101001" => rgb <= "111111";
				  when "11010101101010" => rgb <= "111111";
				  when "11010101101011" => rgb <= "111111";
				  when "11010101101100" => rgb <= "111111";
				  when "11010101101101" => rgb <= "111111";
				  when "11010101101110" => rgb <= "111111";
				  when "11010101101111" => rgb <= "111111";
				  when "11010101110000" => rgb <= "111111";
				  when "11010101110001" => rgb <= "111111";
				  when "11010101110010" => rgb <= "111111";
				  when "11010101110011" => rgb <= "111111";
				  when "11010101110100" => rgb <= "111111";
				  when "11010101110101" => rgb <= "111111";
				  when "11010101110110" => rgb <= "111111";
				  when "11010101110111" => rgb <= "111111";
				  when "11010101111000" => rgb <= "111111";
				  when "11010101111001" => rgb <= "111111";
				  when "11010101111010" => rgb <= "111111";
				  when "11010101111011" => rgb <= "111111";
				  when "11010101111100" => rgb <= "111111";
				  when "11010101111101" => rgb <= "111111";
				  when "11010101111110" => rgb <= "111111";
				  when "11010101111111" => rgb <= "111111";
				  when "11010110000000" => rgb <= "111111";
				  when "11010110000001" => rgb <= "111111";
				  when "11010110000010" => rgb <= "111111";
				  when "11010110000011" => rgb <= "111111";
				  when "11010110000100" => rgb <= "111111";
				  when "11010110000101" => rgb <= "111111";
				  when "11010110000110" => rgb <= "111111";
				  when "11010110000111" => rgb <= "111111";
				  when "11010110001000" => rgb <= "111111";
				  when "11010110001001" => rgb <= "111111";
				  when "11010110001010" => rgb <= "111111";
				  when "11010110001011" => rgb <= "111111";
				  when "11010110001100" => rgb <= "111111";
				  when "11010110001101" => rgb <= "111111";
				  when "11010110001110" => rgb <= "111111";
				  when "11010110001111" => rgb <= "111111";
				  when "11010110010000" => rgb <= "111111";
				  when "11010110010001" => rgb <= "111111";
				  when "11010110010010" => rgb <= "111111";
				  when "11010110010011" => rgb <= "111111";
				  when "11010110010100" => rgb <= "111111";
				  when "11010110010101" => rgb <= "111111";
				  when "11010110010110" => rgb <= "111111";
				  when "11010110010111" => rgb <= "111111";
				  when "11010110011000" => rgb <= "111111";
				  when "11010110011001" => rgb <= "111111";
				  when "11010110011010" => rgb <= "111111";
				  when "11010110011011" => rgb <= "111111";
				  when "11010110011100" => rgb <= "111111";
				  when "11010110011101" => rgb <= "111111";
				  when "11010110011110" => rgb <= "111111";
				  when "11010110011111" => rgb <= "111111";
				  when "11011100000000" => rgb <= "111000";
				  when "11011100000001" => rgb <= "111000";
				  when "11011100000010" => rgb <= "111000";
				  when "11011100000011" => rgb <= "111000";
				  when "11011100000100" => rgb <= "111000";
				  when "11011100000101" => rgb <= "111000";
				  when "11011100000110" => rgb <= "111000";
				  when "11011100000111" => rgb <= "111000";
				  when "11011100001000" => rgb <= "111000";
				  when "11011100001001" => rgb <= "111000";
				  when "11011100001010" => rgb <= "111000";
				  when "11011100001011" => rgb <= "111000";
				  when "11011100001100" => rgb <= "111000";
				  when "11011100001101" => rgb <= "111000";
				  when "11011100001110" => rgb <= "111000";
				  when "11011100001111" => rgb <= "111000";
				  when "11011100010000" => rgb <= "111000";
				  when "11011100010001" => rgb <= "111000";
				  when "11011100010010" => rgb <= "111000";
				  when "11011100010011" => rgb <= "111000";
				  when "11011100010100" => rgb <= "111000";
				  when "11011100010101" => rgb <= "111000";
				  when "11011100010110" => rgb <= "111000";
				  when "11011100010111" => rgb <= "111000";
				  when "11011100011000" => rgb <= "111000";
				  when "11011100011001" => rgb <= "111000";
				  when "11011100011010" => rgb <= "111000";
				  when "11011100011011" => rgb <= "111000";
				  when "11011100011100" => rgb <= "111000";
				  when "11011100011101" => rgb <= "111000";
				  when "11011100011110" => rgb <= "111000";
				  when "11011100011111" => rgb <= "111000";
				  when "11011100100000" => rgb <= "111000";
				  when "11011100100001" => rgb <= "111000";
				  when "11011100100010" => rgb <= "111000";
				  when "11011100100011" => rgb <= "111000";
				  when "11011100100100" => rgb <= "111000";
				  when "11011100100101" => rgb <= "111000";
				  when "11011100100110" => rgb <= "111000";
				  when "11011100100111" => rgb <= "111000";
				  when "11011100101000" => rgb <= "111000";
				  when "11011100101001" => rgb <= "111000";
				  when "11011100101010" => rgb <= "111000";
				  when "11011100101011" => rgb <= "111000";
				  when "11011100101100" => rgb <= "111000";
				  when "11011100101101" => rgb <= "111000";
				  when "11011100101110" => rgb <= "111000";
				  when "11011100101111" => rgb <= "111000";
				  when "11011100110000" => rgb <= "111000";
				  when "11011100110001" => rgb <= "111000";
				  when "11011100110010" => rgb <= "111000";
				  when "11011100110011" => rgb <= "111000";
				  when "11011100110100" => rgb <= "111000";
				  when "11011100110101" => rgb <= "111000";
				  when "11011100110110" => rgb <= "111000";
				  when "11011100110111" => rgb <= "111000";
				  when "11011100111000" => rgb <= "111000";
				  when "11011100111001" => rgb <= "111000";
				  when "11011100111010" => rgb <= "111000";
				  when "11011100111011" => rgb <= "111000";
				  when "11011100111100" => rgb <= "111000";
				  when "11011100111101" => rgb <= "111000";
				  when "11011100111110" => rgb <= "111000";
				  when "11011100111111" => rgb <= "111000";
				  when "11011101000000" => rgb <= "111000";
				  when "11011101000001" => rgb <= "111000";
				  when "11011101000010" => rgb <= "111000";
				  when "11011101000011" => rgb <= "111000";
				  when "11011101000100" => rgb <= "111000";
				  when "11011101000101" => rgb <= "111000";
				  when "11011101000110" => rgb <= "111000";
				  when "11011101000111" => rgb <= "111000";
				  when "11011101001000" => rgb <= "111000";
				  when "11011101001001" => rgb <= "111000";
				  when "11011101001010" => rgb <= "111000";
				  when "11011101001011" => rgb <= "111000";
				  when "11011101001100" => rgb <= "111000";
				  when "11011101001101" => rgb <= "111000";
				  when "11011101001110" => rgb <= "111000";
				  when "11011101001111" => rgb <= "111000";
				  when "11011101010000" => rgb <= "111000";
				  when "11011101010001" => rgb <= "111000";
				  when "11011101010010" => rgb <= "111000";
				  when "11011101010011" => rgb <= "111000";
				  when "11011101010100" => rgb <= "111000";
				  when "11011101010101" => rgb <= "111000";
				  when "11011101010110" => rgb <= "111000";
				  when "11011101010111" => rgb <= "111000";
				  when "11011101011000" => rgb <= "111000";
				  when "11011101011001" => rgb <= "111000";
				  when "11011101011010" => rgb <= "111000";
				  when "11011101011011" => rgb <= "111000";
				  when "11011101011100" => rgb <= "111000";
				  when "11011101011101" => rgb <= "111000";
				  when "11011101011110" => rgb <= "111000";
				  when "11011101011111" => rgb <= "111000";
				  when "11011101100000" => rgb <= "111000";
				  when "11011101100001" => rgb <= "111000";
				  when "11011101100010" => rgb <= "111000";
				  when "11011101100011" => rgb <= "111000";
				  when "11011101100100" => rgb <= "111000";
				  when "11011101100101" => rgb <= "111000";
				  when "11011101100110" => rgb <= "111000";
				  when "11011101100111" => rgb <= "111000";
				  when "11011101101000" => rgb <= "111000";
				  when "11011101101001" => rgb <= "111000";
				  when "11011101101010" => rgb <= "111000";
				  when "11011101101011" => rgb <= "111000";
				  when "11011101101100" => rgb <= "111000";
				  when "11011101101101" => rgb <= "111000";
				  when "11011101101110" => rgb <= "111000";
				  when "11011101101111" => rgb <= "111000";
				  when "11011101110000" => rgb <= "111000";
				  when "11011101110001" => rgb <= "111000";
				  when "11011101110010" => rgb <= "111000";
				  when "11011101110011" => rgb <= "111000";
				  when "11011101110100" => rgb <= "111000";
				  when "11011101110101" => rgb <= "111000";
				  when "11011101110110" => rgb <= "111000";
				  when "11011101110111" => rgb <= "111000";
				  when "11011101111000" => rgb <= "111000";
				  when "11011101111001" => rgb <= "111000";
				  when "11011101111010" => rgb <= "111000";
				  when "11011101111011" => rgb <= "111000";
				  when "11011101111100" => rgb <= "111000";
				  when "11011101111101" => rgb <= "111000";
				  when "11011101111110" => rgb <= "111000";
				  when "11011101111111" => rgb <= "111000";
				  when "11011110000000" => rgb <= "111000";
				  when "11011110000001" => rgb <= "111000";
				  when "11011110000010" => rgb <= "111000";
				  when "11011110000011" => rgb <= "111000";
				  when "11011110000100" => rgb <= "111000";
				  when "11011110000101" => rgb <= "111000";
				  when "11011110000110" => rgb <= "111000";
				  when "11011110000111" => rgb <= "111000";
				  when "11011110001000" => rgb <= "111000";
				  when "11011110001001" => rgb <= "111000";
				  when "11011110001010" => rgb <= "111000";
				  when "11011110001011" => rgb <= "111000";
				  when "11011110001100" => rgb <= "111000";
				  when "11011110001101" => rgb <= "111000";
				  when "11011110001110" => rgb <= "111000";
				  when "11011110001111" => rgb <= "111000";
				  when "11011110010000" => rgb <= "111000";
				  when "11011110010001" => rgb <= "111000";
				  when "11011110010010" => rgb <= "111000";
				  when "11011110010011" => rgb <= "111000";
				  when "11011110010100" => rgb <= "111000";
				  when "11011110010101" => rgb <= "111000";
				  when "11011110010110" => rgb <= "111000";
				  when "11011110010111" => rgb <= "111000";
				  when "11011110011000" => rgb <= "111000";
				  when "11011110011001" => rgb <= "111000";
				  when "11011110011010" => rgb <= "111000";
				  when "11011110011011" => rgb <= "111000";
				  when "11011110011100" => rgb <= "111000";
				  when "11011110011101" => rgb <= "111000";
				  when "11011110011110" => rgb <= "111000";
				  when "11011110011111" => rgb <= "111000";
				  when "11100100000000" => rgb <= "111111";
				  when "11100100000001" => rgb <= "111111";
				  when "11100100000010" => rgb <= "111111";
				  when "11100100000011" => rgb <= "111111";
				  when "11100100000100" => rgb <= "111111";
				  when "11100100000101" => rgb <= "111111";
				  when "11100100000110" => rgb <= "111111";
				  when "11100100000111" => rgb <= "111111";
				  when "11100100001000" => rgb <= "111111";
				  when "11100100001001" => rgb <= "111111";
				  when "11100100001010" => rgb <= "111111";
				  when "11100100001011" => rgb <= "111111";
				  when "11100100001100" => rgb <= "111111";
				  when "11100100001101" => rgb <= "111111";
				  when "11100100001110" => rgb <= "111111";
				  when "11100100001111" => rgb <= "111111";
				  when "11100100010000" => rgb <= "111111";
				  when "11100100010001" => rgb <= "111111";
				  when "11100100010010" => rgb <= "111111";
				  when "11100100010011" => rgb <= "111111";
				  when "11100100010100" => rgb <= "111111";
				  when "11100100010101" => rgb <= "111111";
				  when "11100100010110" => rgb <= "111111";
				  when "11100100010111" => rgb <= "111111";
				  when "11100100011000" => rgb <= "111111";
				  when "11100100011001" => rgb <= "111111";
				  when "11100100011010" => rgb <= "111111";
				  when "11100100011011" => rgb <= "111111";
				  when "11100100011100" => rgb <= "111111";
				  when "11100100011101" => rgb <= "111111";
				  when "11100100011110" => rgb <= "111111";
				  when "11100100011111" => rgb <= "111111";
				  when "11100100100000" => rgb <= "111111";
				  when "11100100100001" => rgb <= "111111";
				  when "11100100100010" => rgb <= "111111";
				  when "11100100100011" => rgb <= "111111";
				  when "11100100100100" => rgb <= "111111";
				  when "11100100100101" => rgb <= "111111";
				  when "11100100100110" => rgb <= "111111";
				  when "11100100100111" => rgb <= "111111";
				  when "11100100101000" => rgb <= "111111";
				  when "11100100101001" => rgb <= "111111";
				  when "11100100101010" => rgb <= "111111";
				  when "11100100101011" => rgb <= "111111";
				  when "11100100101100" => rgb <= "111111";
				  when "11100100101101" => rgb <= "111111";
				  when "11100100101110" => rgb <= "111111";
				  when "11100100101111" => rgb <= "111111";
				  when "11100100110000" => rgb <= "111111";
				  when "11100100110001" => rgb <= "111111";
				  when "11100100110010" => rgb <= "111111";
				  when "11100100110011" => rgb <= "111111";
				  when "11100100110100" => rgb <= "111111";
				  when "11100100110101" => rgb <= "111111";
				  when "11100100110110" => rgb <= "111111";
				  when "11100100110111" => rgb <= "111111";
				  when "11100100111000" => rgb <= "111111";
				  when "11100100111001" => rgb <= "111111";
				  when "11100100111010" => rgb <= "111111";
				  when "11100100111011" => rgb <= "111111";
				  when "11100100111100" => rgb <= "111111";
				  when "11100100111101" => rgb <= "111111";
				  when "11100100111110" => rgb <= "111111";
				  when "11100100111111" => rgb <= "111111";
				  when "11100101000000" => rgb <= "111111";
				  when "11100101000001" => rgb <= "111111";
				  when "11100101000010" => rgb <= "111111";
				  when "11100101000011" => rgb <= "111111";
				  when "11100101000100" => rgb <= "111111";
				  when "11100101000101" => rgb <= "111111";
				  when "11100101000110" => rgb <= "111111";
				  when "11100101000111" => rgb <= "111111";
				  when "11100101001000" => rgb <= "111111";
				  when "11100101001001" => rgb <= "111111";
				  when "11100101001010" => rgb <= "111111";
				  when "11100101001011" => rgb <= "111111";
				  when "11100101001100" => rgb <= "111111";
				  when "11100101001101" => rgb <= "111111";
				  when "11100101001110" => rgb <= "111111";
				  when "11100101001111" => rgb <= "111111";
				  when "11100101010000" => rgb <= "111111";
				  when "11100101010001" => rgb <= "111111";
				  when "11100101010010" => rgb <= "111111";
				  when "11100101010011" => rgb <= "111111";
				  when "11100101010100" => rgb <= "111111";
				  when "11100101010101" => rgb <= "111111";
				  when "11100101010110" => rgb <= "111111";
				  when "11100101010111" => rgb <= "111111";
				  when "11100101011000" => rgb <= "111111";
				  when "11100101011001" => rgb <= "111111";
				  when "11100101011010" => rgb <= "111111";
				  when "11100101011011" => rgb <= "111111";
				  when "11100101011100" => rgb <= "111111";
				  when "11100101011101" => rgb <= "111111";
				  when "11100101011110" => rgb <= "111111";
				  when "11100101011111" => rgb <= "111111";
				  when "11100101100000" => rgb <= "111111";
				  when "11100101100001" => rgb <= "111111";
				  when "11100101100010" => rgb <= "111111";
				  when "11100101100011" => rgb <= "111111";
				  when "11100101100100" => rgb <= "111111";
				  when "11100101100101" => rgb <= "111111";
				  when "11100101100110" => rgb <= "111111";
				  when "11100101100111" => rgb <= "111111";
				  when "11100101101000" => rgb <= "111111";
				  when "11100101101001" => rgb <= "111111";
				  when "11100101101010" => rgb <= "111111";
				  when "11100101101011" => rgb <= "111111";
				  when "11100101101100" => rgb <= "111111";
				  when "11100101101101" => rgb <= "111111";
				  when "11100101101110" => rgb <= "111111";
				  when "11100101101111" => rgb <= "111111";
				  when "11100101110000" => rgb <= "111111";
				  when "11100101110001" => rgb <= "111111";
				  when "11100101110010" => rgb <= "111111";
				  when "11100101110011" => rgb <= "111111";
				  when "11100101110100" => rgb <= "111111";
				  when "11100101110101" => rgb <= "111111";
				  when "11100101110110" => rgb <= "111111";
				  when "11100101110111" => rgb <= "111111";
				  when "11100101111000" => rgb <= "111111";
				  when "11100101111001" => rgb <= "111111";
				  when "11100101111010" => rgb <= "111111";
				  when "11100101111011" => rgb <= "111111";
				  when "11100101111100" => rgb <= "111111";
				  when "11100101111101" => rgb <= "111111";
				  when "11100101111110" => rgb <= "111111";
				  when "11100101111111" => rgb <= "111111";
				  when "11100110000000" => rgb <= "111111";
				  when "11100110000001" => rgb <= "111111";
				  when "11100110000010" => rgb <= "111111";
				  when "11100110000011" => rgb <= "111111";
				  when "11100110000100" => rgb <= "111111";
				  when "11100110000101" => rgb <= "111111";
				  when "11100110000110" => rgb <= "111111";
				  when "11100110000111" => rgb <= "111111";
				  when "11100110001000" => rgb <= "111111";
				  when "11100110001001" => rgb <= "111111";
				  when "11100110001010" => rgb <= "111111";
				  when "11100110001011" => rgb <= "111111";
				  when "11100110001100" => rgb <= "111111";
				  when "11100110001101" => rgb <= "111111";
				  when "11100110001110" => rgb <= "111111";
				  when "11100110001111" => rgb <= "111111";
				  when "11100110010000" => rgb <= "111111";
				  when "11100110010001" => rgb <= "111111";
				  when "11100110010010" => rgb <= "111111";
				  when "11100110010011" => rgb <= "111111";
				  when "11100110010100" => rgb <= "111111";
				  when "11100110010101" => rgb <= "111111";
				  when "11100110010110" => rgb <= "111111";
				  when "11100110010111" => rgb <= "111111";
				  when "11100110011000" => rgb <= "111111";
				  when "11100110011001" => rgb <= "111111";
				  when "11100110011010" => rgb <= "111111";
				  when "11100110011011" => rgb <= "111111";
				  when "11100110011100" => rgb <= "111111";
				  when "11100110011101" => rgb <= "111111";
				  when "11100110011110" => rgb <= "111111";
				  when "11100110011111" => rgb <= "111111";
				  when "11101000000000" => rgb <= "111111";
				  when "11101000000001" => rgb <= "111111";
				  when "11101000000010" => rgb <= "111111";
				  when "11101000000011" => rgb <= "111111";
				  when "11101000000100" => rgb <= "111111";
				  when "11101000000101" => rgb <= "111111";
				  when "11101000000110" => rgb <= "111111";
				  when "11101000000111" => rgb <= "111111";
				  when "11101000001000" => rgb <= "111111";
				  when "11101000001001" => rgb <= "111111";
				  when "11101000001010" => rgb <= "111111";
				  when "11101000001011" => rgb <= "111111";
				  when "11101000001100" => rgb <= "111111";
				  when "11101000001101" => rgb <= "111111";
				  when "11101000001110" => rgb <= "111111";
				  when "11101000001111" => rgb <= "111111";
				  when "11101000010000" => rgb <= "111111";
				  when "11101000010001" => rgb <= "111111";
				  when "11101000010010" => rgb <= "111111";
				  when "11101000010011" => rgb <= "111111";
				  when "11101000010100" => rgb <= "111111";
				  when "11101000010101" => rgb <= "111111";
				  when "11101000010110" => rgb <= "111111";
				  when "11101000010111" => rgb <= "111111";
				  when "11101000011000" => rgb <= "111111";
				  when "11101000011001" => rgb <= "111111";
				  when "11101000011010" => rgb <= "111111";
				  when "11101000011011" => rgb <= "111111";
				  when "11101000011100" => rgb <= "111111";
				  when "11101000011101" => rgb <= "111111";
				  when "11101000011110" => rgb <= "111111";
				  when "11101000011111" => rgb <= "111111";
				  when "11101000100000" => rgb <= "111111";
				  when "11101000100001" => rgb <= "111111";
				  when "11101000100010" => rgb <= "111111";
				  when "11101000100011" => rgb <= "111111";
				  when "11101000100100" => rgb <= "111111";
				  when "11101000100101" => rgb <= "111111";
				  when "11101000100110" => rgb <= "111111";
				  when "11101000100111" => rgb <= "111111";
				  when "11101000101000" => rgb <= "111111";
				  when "11101000101001" => rgb <= "111111";
				  when "11101000101010" => rgb <= "111111";
				  when "11101000101011" => rgb <= "111111";
				  when "11101000101100" => rgb <= "111111";
				  when "11101000101101" => rgb <= "111111";
				  when "11101000101110" => rgb <= "111111";
				  when "11101000101111" => rgb <= "111111";
				  when "11101000110000" => rgb <= "111111";
				  when "11101000110001" => rgb <= "111111";
				  when "11101000110010" => rgb <= "111111";
				  when "11101000110011" => rgb <= "111111";
				  when "11101000110100" => rgb <= "111111";
				  when "11101000110101" => rgb <= "111111";
				  when "11101000110110" => rgb <= "111111";
				  when "11101000110111" => rgb <= "111111";
				  when "11101000111000" => rgb <= "111111";
				  when "11101000111001" => rgb <= "111111";
				  when "11101000111010" => rgb <= "111111";
				  when "11101000111011" => rgb <= "111111";
				  when "11101000111100" => rgb <= "111111";
				  when "11101000111101" => rgb <= "111111";
				  when "11101000111110" => rgb <= "111111";
				  when "11101000111111" => rgb <= "111111";
				  when "11101001000000" => rgb <= "111111";
				  when "11101001000001" => rgb <= "111111";
				  when "11101001000010" => rgb <= "111111";
				  when "11101001000011" => rgb <= "111111";
				  when "11101001000100" => rgb <= "111111";
				  when "11101001000101" => rgb <= "111111";
				  when "11101001000110" => rgb <= "111111";
				  when "11101001000111" => rgb <= "111111";
				  when "11101001001000" => rgb <= "111111";
				  when "11101001001001" => rgb <= "111111";
				  when "11101001001010" => rgb <= "111111";
				  when "11101001001011" => rgb <= "111111";
				  when "11101001001100" => rgb <= "111111";
				  when "11101001001101" => rgb <= "111111";
				  when "11101001001110" => rgb <= "111111";
				  when "11101001001111" => rgb <= "111111";
				  when "11101001010000" => rgb <= "111111";
				  when "11101001010001" => rgb <= "111111";
				  when "11101001010010" => rgb <= "111111";
				  when "11101001010011" => rgb <= "111111";
				  when "11101001010100" => rgb <= "111111";
				  when "11101001010101" => rgb <= "111111";
				  when "11101001010110" => rgb <= "111111";
				  when "11101001010111" => rgb <= "111111";
				  when "11101001011000" => rgb <= "111111";
				  when "11101001011001" => rgb <= "111111";
				  when "11101001011010" => rgb <= "111111";
				  when "11101001011011" => rgb <= "111111";
				  when "11101001011100" => rgb <= "111111";
				  when "11101001011101" => rgb <= "111111";
				  when "11101001011110" => rgb <= "111111";
				  when "11101001011111" => rgb <= "111111";
				  when "11101001100000" => rgb <= "111111";
				  when "11101001100001" => rgb <= "111111";
				  when "11101001100010" => rgb <= "111111";
				  when "11101001100011" => rgb <= "111111";
				  when "11101001100100" => rgb <= "111111";
				  when "11101001100101" => rgb <= "111111";
				  when "11101001100110" => rgb <= "111111";
				  when "11101001100111" => rgb <= "111111";
				  when "11101001101000" => rgb <= "111111";
				  when "11101001101001" => rgb <= "111111";
				  when "11101001101010" => rgb <= "111111";
				  when "11101001101011" => rgb <= "111111";
				  when "11101001101100" => rgb <= "111111";
				  when "11101001101101" => rgb <= "111111";
				  when "11101001101110" => rgb <= "111111";
				  when "11101001101111" => rgb <= "111111";
				  when "11101001110000" => rgb <= "111111";
				  when "11101001110001" => rgb <= "111111";
				  when "11101001110010" => rgb <= "111111";
				  when "11101001110011" => rgb <= "111111";
				  when "11101001110100" => rgb <= "111111";
				  when "11101001110101" => rgb <= "111111";
				  when "11101001110110" => rgb <= "111111";
				  when "11101001110111" => rgb <= "111111";
				  when "11101001111000" => rgb <= "111111";
				  when "11101001111001" => rgb <= "111111";
				  when "11101001111010" => rgb <= "111111";
				  when "11101001111011" => rgb <= "111111";
				  when "11101001111100" => rgb <= "111111";
				  when "11101001111101" => rgb <= "111111";
				  when "11101001111110" => rgb <= "111111";
				  when "11101001111111" => rgb <= "111111";
				  when "11101010000000" => rgb <= "111111";
				  when "11101010000001" => rgb <= "111111";
				  when "11101010000010" => rgb <= "111111";
				  when "11101010000011" => rgb <= "111111";
				  when "11101010000100" => rgb <= "111111";
				  when "11101010000101" => rgb <= "111111";
				  when "11101010000110" => rgb <= "111111";
				  when "11101010000111" => rgb <= "111111";
				  when "11101010001000" => rgb <= "111111";
				  when "11101010001001" => rgb <= "111111";
				  when "11101010001010" => rgb <= "111111";
				  when "11101010001011" => rgb <= "111111";
				  when "11101010001100" => rgb <= "111111";
				  when "11101010001101" => rgb <= "111111";
				  when "11101010001110" => rgb <= "111111";
				  when "11101010001111" => rgb <= "111111";
				  when "11101010010000" => rgb <= "111111";
				  when "11101010010001" => rgb <= "111111";
				  when "11101010010010" => rgb <= "111111";
				  when "11101010010011" => rgb <= "111111";
				  when "11101010010100" => rgb <= "111111";
				  when "11101010010101" => rgb <= "111111";
				  when "11101010010110" => rgb <= "111111";
				  when "11101010010111" => rgb <= "111111";
				  when "11101010011000" => rgb <= "111111";
				  when "11101010011001" => rgb <= "111111";
				  when "11101010011010" => rgb <= "111111";
				  when "11101010011011" => rgb <= "111111";
				  when "11101010011100" => rgb <= "111111";
				  when "11101010011101" => rgb <= "111111";
				  when "11101010011110" => rgb <= "111111";
				  when "11101010011111" => rgb <= "111111";
				  when "11101100000000" => rgb <= "111111";
				  when "11101100000001" => rgb <= "111111";
				  when "11101100000010" => rgb <= "111111";
				  when "11101100000011" => rgb <= "111111";
				  when "11101100000100" => rgb <= "111111";
				  when "11101100000101" => rgb <= "111111";
				  when "11101100000110" => rgb <= "111111";
				  when "11101100000111" => rgb <= "111111";
				  when "11101100001000" => rgb <= "111111";
				  when "11101100001001" => rgb <= "111111";
				  when "11101100001010" => rgb <= "111111";
				  when "11101100001011" => rgb <= "111111";
				  when "11101100001100" => rgb <= "111111";
				  when "11101100001101" => rgb <= "111111";
				  when "11101100001110" => rgb <= "111111";
				  when "11101100001111" => rgb <= "111111";
				  when "11101100010000" => rgb <= "111111";
				  when "11101100010001" => rgb <= "111111";
				  when "11101100010010" => rgb <= "111111";
				  when "11101100010011" => rgb <= "111111";
				  when "11101100010100" => rgb <= "111111";
				  when "11101100010101" => rgb <= "111111";
				  when "11101100010110" => rgb <= "111111";
				  when "11101100010111" => rgb <= "111111";
				  when "11101100011000" => rgb <= "111111";
				  when "11101100011001" => rgb <= "111111";
				  when "11101100011010" => rgb <= "111111";
				  when "11101100011011" => rgb <= "111111";
				  when "11101100011100" => rgb <= "111111";
				  when "11101100011101" => rgb <= "111111";
				  when "11101100011110" => rgb <= "111111";
				  when "11101100011111" => rgb <= "111111";
				  when "11101100100000" => rgb <= "111111";
				  when "11101100100001" => rgb <= "111111";
				  when "11101100100010" => rgb <= "111111";
				  when "11101100100011" => rgb <= "111111";
				  when "11101100100100" => rgb <= "111111";
				  when "11101100100101" => rgb <= "111111";
				  when "11101100100110" => rgb <= "111111";
				  when "11101100100111" => rgb <= "111111";
				  when "11101100101000" => rgb <= "111111";
				  when "11101100101001" => rgb <= "111111";
				  when "11101100101010" => rgb <= "111111";
				  when "11101100101011" => rgb <= "111111";
				  when "11101100101100" => rgb <= "111111";
				  when "11101100101101" => rgb <= "111111";
				  when "11101100101110" => rgb <= "111111";
				  when "11101100101111" => rgb <= "111111";
				  when "11101100110000" => rgb <= "111111";
				  when "11101100110001" => rgb <= "111111";
				  when "11101100110010" => rgb <= "111111";
				  when "11101100110011" => rgb <= "111111";
				  when "11101100110100" => rgb <= "111111";
				  when "11101100110101" => rgb <= "111111";
				  when "11101100110110" => rgb <= "111111";
				  when "11101100110111" => rgb <= "111111";
				  when "11101100111000" => rgb <= "111111";
				  when "11101100111001" => rgb <= "111111";
				  when "11101100111010" => rgb <= "111111";
				  when "11101100111011" => rgb <= "111111";
				  when "11101100111100" => rgb <= "111111";
				  when "11101100111101" => rgb <= "111111";
				  when "11101100111110" => rgb <= "111111";
				  when "11101100111111" => rgb <= "111111";
				  when "11101101000000" => rgb <= "111111";
				  when "11101101000001" => rgb <= "111111";
				  when "11101101000010" => rgb <= "111111";
				  when "11101101000011" => rgb <= "111111";
				  when "11101101000100" => rgb <= "111111";
				  when "11101101000101" => rgb <= "111111";
				  when "11101101000110" => rgb <= "111111";
				  when "11101101000111" => rgb <= "111111";
				  when "11101101001000" => rgb <= "111111";
				  when "11101101001001" => rgb <= "111111";
				  when "11101101001010" => rgb <= "111111";
				  when "11101101001011" => rgb <= "111111";
				  when "11101101001100" => rgb <= "111111";
				  when "11101101001101" => rgb <= "111111";
				  when "11101101001110" => rgb <= "111111";
				  when "11101101001111" => rgb <= "111111";
				  when "11101101010000" => rgb <= "111111";
				  when "11101101010001" => rgb <= "111111";
				  when "11101101010010" => rgb <= "111111";
				  when "11101101010011" => rgb <= "111111";
				  when "11101101010100" => rgb <= "111111";
				  when "11101101010101" => rgb <= "111111";
				  when "11101101010110" => rgb <= "111111";
				  when "11101101010111" => rgb <= "111111";
				  when "11101101011000" => rgb <= "111111";
				  when "11101101011001" => rgb <= "111111";
				  when "11101101011010" => rgb <= "111111";
				  when "11101101011011" => rgb <= "111111";
				  when "11101101011100" => rgb <= "111111";
				  when "11101101011101" => rgb <= "111111";
				  when "11101101011110" => rgb <= "111111";
				  when "11101101011111" => rgb <= "111111";
				  when "11101101100000" => rgb <= "111111";
				  when "11101101100001" => rgb <= "111111";
				  when "11101101100010" => rgb <= "111111";
				  when "11101101100011" => rgb <= "111111";
				  when "11101101100100" => rgb <= "111111";
				  when "11101101100101" => rgb <= "111111";
				  when "11101101100110" => rgb <= "111111";
				  when "11101101100111" => rgb <= "111111";
				  when "11101101101000" => rgb <= "111111";
				  when "11101101101001" => rgb <= "111111";
				  when "11101101101010" => rgb <= "111111";
				  when "11101101101011" => rgb <= "111111";
				  when "11101101101100" => rgb <= "111111";
				  when "11101101101101" => rgb <= "111111";
				  when "11101101101110" => rgb <= "111111";
				  when "11101101101111" => rgb <= "111111";
				  when "11101101110000" => rgb <= "111111";
				  when "11101101110001" => rgb <= "111111";
				  when "11101101110010" => rgb <= "111111";
				  when "11101101110011" => rgb <= "111111";
				  when "11101101110100" => rgb <= "111111";
				  when "11101101110101" => rgb <= "111111";
				  when "11101101110110" => rgb <= "111111";
				  when "11101101110111" => rgb <= "111111";
				  when "11101101111000" => rgb <= "111111";
				  when "11101101111001" => rgb <= "111111";
				  when "11101101111010" => rgb <= "111111";
				  when "11101101111011" => rgb <= "111111";
				  when "11101101111100" => rgb <= "111111";
				  when "11101101111101" => rgb <= "111111";
				  when "11101101111110" => rgb <= "111111";
				  when "11101101111111" => rgb <= "111111";
				  when "11101110000000" => rgb <= "111111";
				  when "11101110000001" => rgb <= "111111";
				  when "11101110000010" => rgb <= "111111";
				  when "11101110000011" => rgb <= "111111";
				  when "11101110000100" => rgb <= "111111";
				  when "11101110000101" => rgb <= "111111";
				  when "11101110000110" => rgb <= "111111";
				  when "11101110000111" => rgb <= "111111";
				  when "11101110001000" => rgb <= "111111";
				  when "11101110001001" => rgb <= "111111";
				  when "11101110001010" => rgb <= "111111";
				  when "11101110001011" => rgb <= "111111";
				  when "11101110001100" => rgb <= "111111";
				  when "11101110001101" => rgb <= "111111";
				  when "11101110001110" => rgb <= "111111";
				  when "11101110001111" => rgb <= "111111";
				  when "11101110010000" => rgb <= "111111";
				  when "11101110010001" => rgb <= "111111";
				  when "11101110010010" => rgb <= "111111";
				  when "11101110010011" => rgb <= "111111";
				  when "11101110010100" => rgb <= "111111";
				  when "11101110010101" => rgb <= "111111";
				  when "11101110010110" => rgb <= "111111";
				  when "11101110010111" => rgb <= "111111";
				  when "11101110011000" => rgb <= "111111";
				  when "11101110011001" => rgb <= "111111";
				  when "11101110011010" => rgb <= "111111";
				  when "11101110011011" => rgb <= "111111";
				  when "11101110011100" => rgb <= "111111";
				  when "11101110011101" => rgb <= "111111";
				  when "11101110011110" => rgb <= "111111";
				  when "11101110011111" => rgb <= "111111";
				  when others => rgb <= "000000";
			end case;
		end if;
	end process;
	location <= std_logic_vector(col_idx) & std_logic_vector(row_idx);
end;
