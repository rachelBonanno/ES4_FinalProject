library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity gameoverp1_rom is
  port(
	  clk : in std_logic;
	  row_idx: in unsigned(6 downto 0);
	  col_idx : in unsigned(5 downto 0); 
	  rgb : out std_logic_vector(5 downto 0)
	  );
end gameoverp1_rom;

architecture synth of gameoverp1_rom is

signal location : std_logic_vector(12 downto 0);
begin
	process (clk) begin
		if rising_edge(clk) then
			case location is
				                when "0010000000110" => rgb <= "100001";
                when "0010000000111" => rgb <= "100100";
                when "0010000001000" => rgb <= "100100";
                when "0010000001001" => rgb <= "100100";
                when "0010000001010" => rgb <= "100100";
                when "0010000001011" => rgb <= "100001";
                when "0010000001100" => rgb <= "100001";
                when "0010000001101" => rgb <= "100001";
                when "0010000001110" => rgb <= "100001";
                when "0010000001111" => rgb <= "010000";
                when "0010000010000" => rgb <= "100001";
                when "0010000010001" => rgb <= "100001";
                when "0010000010110" => rgb <= "100001";
                when "0010000010111" => rgb <= "100001";
                when "0010000011000" => rgb <= "100001";
                when "0010000011001" => rgb <= "100100";
                when "0010000011110" => rgb <= "100001";
                when "0010000011111" => rgb <= "100001";
                when "0010000100000" => rgb <= "100001";
                when "0010000100001" => rgb <= "100001";
                when "0010000100110" => rgb <= "100001";
                when "0010000100111" => rgb <= "100001";
                when "0010000101000" => rgb <= "100001";
                when "0010000101001" => rgb <= "100001";
                when "0010000101010" => rgb <= "010000";
                when "0010000101011" => rgb <= "010000";
                when "0010000101100" => rgb <= "100001";
                when "0010000101101" => rgb <= "100001";
                when "0010000110010" => rgb <= "100001";
                when "0010000110011" => rgb <= "100001";
                when "0010000110100" => rgb <= "100001";
                when "0010000110101" => rgb <= "100001";
                when "0010000111010" => rgb <= "100001";
                when "0010000111011" => rgb <= "100001";
                when "0010000111100" => rgb <= "100001";
                when "0010000111101" => rgb <= "100001";
                when "0010001000010" => rgb <= "100001";
                when "0010001000011" => rgb <= "100001";
                when "0010001000100" => rgb <= "100001";
                when "0010001000101" => rgb <= "100001";
                when "0010001000110" => rgb <= "100001";
                when "0010001000111" => rgb <= "100001";
                when "0010001001000" => rgb <= "100100";
                when "0010001001001" => rgb <= "100100";
                when "0010010000110" => rgb <= "010000";
                when "0010010000111" => rgb <= "010000";
                when "0010010001000" => rgb <= "100001";
                when "0010010001001" => rgb <= "100001";
                when "0010010001010" => rgb <= "100001";
                when "0010010001011" => rgb <= "100001";
                when "0010010001100" => rgb <= "100001";
                when "0010010001101" => rgb <= "100001";
                when "0010010001110" => rgb <= "100001";
                when "0010010001111" => rgb <= "100001";
                when "0010010010000" => rgb <= "100001";
                when "0010010010001" => rgb <= "100001";
                when "0010010010110" => rgb <= "100001";
                when "0010010010111" => rgb <= "100001";
                when "0010010011000" => rgb <= "100001";
                when "0010010011001" => rgb <= "100001";
                when "0010010011110" => rgb <= "100001";
                when "0010010011111" => rgb <= "100001";
                when "0010010100000" => rgb <= "100001";
                when "0010010100001" => rgb <= "100001";
                when "0010010100110" => rgb <= "100001";
                when "0010010100111" => rgb <= "100100";
                when "0010010101000" => rgb <= "100100";
                when "0010010101001" => rgb <= "100100";
                when "0010010101010" => rgb <= "100100";
                when "0010010101011" => rgb <= "100001";
                when "0010010101100" => rgb <= "100001";
                when "0010010101101" => rgb <= "100001";
                when "0010010110010" => rgb <= "100001";
                when "0010010110011" => rgb <= "100100";
                when "0010010110100" => rgb <= "100100";
                when "0010010110101" => rgb <= "100001";
                when "0010010111001" => rgb <= "100001";
                when "0010010111010" => rgb <= "100100";
                when "0010010111011" => rgb <= "100001";
                when "0010010111100" => rgb <= "010000";
                when "0010010111101" => rgb <= "100001";
                when "0010011000010" => rgb <= "100100";
                when "0010011000011" => rgb <= "100001";
                when "0010011000100" => rgb <= "100001";
                when "0010011000101" => rgb <= "100001";
                when "0010011000110" => rgb <= "100100";
                when "0010011000111" => rgb <= "100100";
                when "0010011001000" => rgb <= "100100";
                when "0010011001001" => rgb <= "100001";
                when "0010100000110" => rgb <= "100100";
                when "0010100000111" => rgb <= "100100";
                when "0010100001000" => rgb <= "100100";
                when "0010100001001" => rgb <= "100001";
                when "0010100001010" => rgb <= "100001";
                when "0010100001011" => rgb <= "100001";
                when "0010100001100" => rgb <= "100001";
                when "0010100001101" => rgb <= "100100";
                when "0010100001110" => rgb <= "100100";
                when "0010100001111" => rgb <= "100100";
                when "0010100010000" => rgb <= "100100";
                when "0010100010001" => rgb <= "100001";
                when "0010100010110" => rgb <= "100001";
                when "0010100010111" => rgb <= "100001";
                when "0010100011000" => rgb <= "100001";
                when "0010100011001" => rgb <= "100001";
                when "0010100011110" => rgb <= "100001";
                when "0010100011111" => rgb <= "010000";
                when "0010100100000" => rgb <= "010000";
                when "0010100100001" => rgb <= "100001";
                when "0010100100110" => rgb <= "100001";
                when "0010100100111" => rgb <= "010000";
                when "0010100101000" => rgb <= "100001";
                when "0010100101001" => rgb <= "100001";
                when "0010100101010" => rgb <= "100001";
                when "0010100101011" => rgb <= "100001";
                when "0010100101100" => rgb <= "100001";
                when "0010100101101" => rgb <= "100001";
                when "0010100110010" => rgb <= "100001";
                when "0010100110011" => rgb <= "100001";
                when "0010100110100" => rgb <= "100100";
                when "0010100110101" => rgb <= "100001";
                when "0010100111000" => rgb <= "100001";
                when "0010100111001" => rgb <= "100001";
                when "0010100111010" => rgb <= "100001";
                when "0010100111011" => rgb <= "100001";
                when "0010100111100" => rgb <= "100001";
                when "0010101000010" => rgb <= "100001";
                when "0010101000011" => rgb <= "100001";
                when "0010101000100" => rgb <= "100001";
                when "0010101000101" => rgb <= "010000";
                when "0010101000110" => rgb <= "010000";
                when "0010101000111" => rgb <= "010000";
                when "0010101001000" => rgb <= "010000";
                when "0010101001001" => rgb <= "100001";
                when "0010110000110" => rgb <= "100001";
                when "0010110000111" => rgb <= "010000";
                when "0010110001000" => rgb <= "100100";
                when "0010110001001" => rgb <= "100100";
                when "0010110001010" => rgb <= "100001";
                when "0010110001011" => rgb <= "100001";
                when "0010110001100" => rgb <= "010000";
                when "0010110001101" => rgb <= "010000";
                when "0010110001110" => rgb <= "100001";
                when "0010110001111" => rgb <= "010000";
                when "0010110010000" => rgb <= "010000";
                when "0010110010001" => rgb <= "100001";
                when "0010110010110" => rgb <= "100001";
                when "0010110010111" => rgb <= "100100";
                when "0010110011000" => rgb <= "100001";
                when "0010110011001" => rgb <= "100001";
                when "0010110011110" => rgb <= "100001";
                when "0010110011111" => rgb <= "100100";
                when "0010110100000" => rgb <= "100001";
                when "0010110100001" => rgb <= "100001";
                when "0010110100110" => rgb <= "100001";
                when "0010110100111" => rgb <= "100001";
                when "0010110101000" => rgb <= "100001";
                when "0010110101001" => rgb <= "100001";
                when "0010110101010" => rgb <= "100001";
                when "0010110101011" => rgb <= "100001";
                when "0010110101100" => rgb <= "100001";
                when "0010110101101" => rgb <= "100001";
                when "0010110110010" => rgb <= "100001";
                when "0010110110011" => rgb <= "100001";
                when "0010110110100" => rgb <= "010000";
                when "0010110110101" => rgb <= "010000";
                when "0010110110111" => rgb <= "100001";
                when "0010110111000" => rgb <= "010000";
                when "0010110111001" => rgb <= "010000";
                when "0010110111010" => rgb <= "100001";
                when "0010110111011" => rgb <= "100001";
                when "0010111000010" => rgb <= "100001";
                when "0010111000011" => rgb <= "100001";
                when "0010111000100" => rgb <= "100001";
                when "0010111000101" => rgb <= "100001";
                when "0010111000110" => rgb <= "100001";
                when "0010111000111" => rgb <= "100001";
                when "0010111001000" => rgb <= "100001";
                when "0010111001001" => rgb <= "100001";
                when "0011000001010" => rgb <= "100001";
                when "0011000001011" => rgb <= "100001";
                when "0011000001100" => rgb <= "100001";
                when "0011000001101" => rgb <= "100001";
                when "0011000010110" => rgb <= "100001";
                when "0011000010111" => rgb <= "100001";
                when "0011000011000" => rgb <= "100001";
                when "0011000011001" => rgb <= "100001";
                when "0011000011110" => rgb <= "100001";
                when "0011000011111" => rgb <= "100001";
                when "0011000100000" => rgb <= "100001";
                when "0011000100001" => rgb <= "100001";
                when "0011000100110" => rgb <= "100100";
                when "0011000100111" => rgb <= "100100";
                when "0011000101000" => rgb <= "100100";
                when "0011000101001" => rgb <= "100001";
                when "0011000110010" => rgb <= "100001";
                when "0011000110011" => rgb <= "010000";
                when "0011000110100" => rgb <= "010000";
                when "0011000110101" => rgb <= "100001";
                when "0011000110110" => rgb <= "100001";
                when "0011000110111" => rgb <= "100100";
                when "0011000111000" => rgb <= "100100";
                when "0011000111001" => rgb <= "100100";
                when "0011000111010" => rgb <= "100001";
                when "0011001000010" => rgb <= "100001";
                when "0011001000011" => rgb <= "100001";
                when "0011001000100" => rgb <= "100100";
                when "0011001000101" => rgb <= "100001";
                when "0011010001010" => rgb <= "100001";
                when "0011010001011" => rgb <= "100001";
                when "0011010001100" => rgb <= "100001";
                when "0011010001101" => rgb <= "100001";
                when "0011010010110" => rgb <= "010000";
                when "0011010010111" => rgb <= "010000";
                when "0011010011000" => rgb <= "100001";
                when "0011010011001" => rgb <= "100001";
                when "0011010011110" => rgb <= "100001";
                when "0011010011111" => rgb <= "100100";
                when "0011010100000" => rgb <= "100001";
                when "0011010100001" => rgb <= "100001";
                when "0011010100110" => rgb <= "100001";
                when "0011010100111" => rgb <= "100001";
                when "0011010101000" => rgb <= "100001";
                when "0011010101001" => rgb <= "100001";
                when "0011010110010" => rgb <= "100001";
                when "0011010110011" => rgb <= "100001";
                when "0011010110100" => rgb <= "100001";
                when "0011010110101" => rgb <= "100001";
                when "0011010110110" => rgb <= "100001";
                when "0011010110111" => rgb <= "100001";
                when "0011010111000" => rgb <= "100001";
                when "0011010111001" => rgb <= "100001";
                when "0011011000010" => rgb <= "100001";
                when "0011011000011" => rgb <= "100001";
                when "0011011000100" => rgb <= "100001";
                when "0011011000101" => rgb <= "100001";
                when "0011100001010" => rgb <= "100001";
                when "0011100001011" => rgb <= "100001";
                when "0011100001100" => rgb <= "100001";
                when "0011100001101" => rgb <= "100001";
                when "0011100010110" => rgb <= "100001";
                when "0011100010111" => rgb <= "100001";
                when "0011100011000" => rgb <= "100001";
                when "0011100011001" => rgb <= "100001";
                when "0011100011110" => rgb <= "100001";
                when "0011100011111" => rgb <= "100001";
                when "0011100100000" => rgb <= "010000";
                when "0011100100001" => rgb <= "100001";
                when "0011100100110" => rgb <= "100001";
                when "0011100100111" => rgb <= "100100";
                when "0011100101000" => rgb <= "100001";
                when "0011100101001" => rgb <= "100001";
                when "0011100101010" => rgb <= "100001";
                when "0011100101011" => rgb <= "010000";
                when "0011100101100" => rgb <= "010000";
                when "0011100101101" => rgb <= "010000";
                when "0011100110010" => rgb <= "100001";
                when "0011100110011" => rgb <= "100001";
                when "0011100110100" => rgb <= "100001";
                when "0011100110101" => rgb <= "100001";
                when "0011100110110" => rgb <= "100001";
                when "0011100110111" => rgb <= "100001";
                when "0011100111000" => rgb <= "100001";
                when "0011101000010" => rgb <= "100001";
                when "0011101000011" => rgb <= "100001";
                when "0011101000100" => rgb <= "100001";
                when "0011101000101" => rgb <= "100001";
                when "0011101000110" => rgb <= "100001";
                when "0011101000111" => rgb <= "100001";
                when "0011101001000" => rgb <= "100001";
                when "0011101001001" => rgb <= "100001";
                when "0011110001010" => rgb <= "100001";
                when "0011110001011" => rgb <= "100001";
                when "0011110001100" => rgb <= "100001";
                when "0011110001101" => rgb <= "100001";
                when "0011110010110" => rgb <= "100001";
                when "0011110010111" => rgb <= "100100";
                when "0011110011000" => rgb <= "100100";
                when "0011110011001" => rgb <= "100001";
                when "0011110011110" => rgb <= "010000";
                when "0011110011111" => rgb <= "010000";
                when "0011110100000" => rgb <= "100001";
                when "0011110100001" => rgb <= "100100";
                when "0011110100110" => rgb <= "100001";
                when "0011110100111" => rgb <= "100001";
                when "0011110101000" => rgb <= "100001";
                when "0011110101001" => rgb <= "100001";
                when "0011110101010" => rgb <= "100100";
                when "0011110101011" => rgb <= "100100";
                when "0011110101100" => rgb <= "100100";
                when "0011110101101" => rgb <= "100001";
                when "0011110110010" => rgb <= "100001";
                when "0011110110011" => rgb <= "100001";
                when "0011110110100" => rgb <= "100001";
                when "0011110110101" => rgb <= "010000";
                when "0011110110110" => rgb <= "010000";
                when "0011110110111" => rgb <= "010000";
                when "0011110111000" => rgb <= "100001";
                when "0011111000010" => rgb <= "100001";
                when "0011111000011" => rgb <= "100001";
                when "0011111000100" => rgb <= "100001";
                when "0011111000101" => rgb <= "100001";
                when "0011111000110" => rgb <= "010000";
                when "0011111000111" => rgb <= "100001";
                when "0011111001000" => rgb <= "100100";
                when "0011111001001" => rgb <= "100100";
                when "0100000001010" => rgb <= "010000";
                when "0100000001011" => rgb <= "100001";
                when "0100000001100" => rgb <= "100001";
                when "0100000001101" => rgb <= "100001";
                when "0100000010110" => rgb <= "100001";
                when "0100000010111" => rgb <= "100001";
                when "0100000011000" => rgb <= "100100";
                when "0100000011001" => rgb <= "100001";
                when "0100000011110" => rgb <= "100001";
                when "0100000011111" => rgb <= "100001";
                when "0100000100000" => rgb <= "100001";
                when "0100000100001" => rgb <= "100001";
                when "0100000101010" => rgb <= "100001";
                when "0100000101011" => rgb <= "100001";
                when "0100000101100" => rgb <= "100100";
                when "0100000101101" => rgb <= "100100";
                when "0100000110010" => rgb <= "100001";
                when "0100000110011" => rgb <= "100100";
                when "0100000110100" => rgb <= "100100";
                when "0100000110101" => rgb <= "100100";
                when "0100000110110" => rgb <= "100100";
                when "0100000110111" => rgb <= "100100";
                when "0100000111000" => rgb <= "100001";
                when "0100000111001" => rgb <= "100001";
                when "0100001000110" => rgb <= "100001";
                when "0100001000111" => rgb <= "100001";
                when "0100001001000" => rgb <= "010000";
                when "0100001001001" => rgb <= "100001";
                when "0100010001010" => rgb <= "100001";
                when "0100010001011" => rgb <= "100001";
                when "0100010001100" => rgb <= "100001";
                when "0100010001101" => rgb <= "100001";
                when "0100010010110" => rgb <= "100001";
                when "0100010010111" => rgb <= "100001";
                when "0100010011000" => rgb <= "100001";
                when "0100010011001" => rgb <= "100001";
                when "0100010011110" => rgb <= "100001";
                when "0100010011111" => rgb <= "100001";
                when "0100010100000" => rgb <= "100001";
                when "0100010100001" => rgb <= "100001";
                when "0100010101010" => rgb <= "010000";
                when "0100010101011" => rgb <= "010000";
                when "0100010101100" => rgb <= "100001";
                when "0100010101101" => rgb <= "100001";
                when "0100010110010" => rgb <= "100001";
                when "0100010110011" => rgb <= "100001";
                when "0100010110100" => rgb <= "100001";
                when "0100010110101" => rgb <= "100001";
                when "0100010110110" => rgb <= "100001";
                when "0100010110111" => rgb <= "100100";
                when "0100010111000" => rgb <= "100100";
                when "0100010111001" => rgb <= "100100";
                when "0100010111010" => rgb <= "010000";
                when "0100011000110" => rgb <= "100001";
                when "0100011000111" => rgb <= "100100";
                when "0100011001000" => rgb <= "100001";
                when "0100011001001" => rgb <= "100001";
                when "0100100001010" => rgb <= "100001";
                when "0100100001011" => rgb <= "100001";
                when "0100100001100" => rgb <= "100001";
                when "0100100001101" => rgb <= "100001";
                when "0100100010110" => rgb <= "100001";
                when "0100100010111" => rgb <= "010000";
                when "0100100011000" => rgb <= "010000";
                when "0100100011001" => rgb <= "100001";
                when "0100100011010" => rgb <= "100001";
                when "0100100011011" => rgb <= "100100";
                when "0100100011100" => rgb <= "100100";
                when "0100100011101" => rgb <= "100100";
                when "0100100011110" => rgb <= "100001";
                when "0100100011111" => rgb <= "010000";
                when "0100100100000" => rgb <= "010000";
                when "0100100100001" => rgb <= "100001";
                when "0100100100110" => rgb <= "100001";
                when "0100100100111" => rgb <= "100100";
                when "0100100101000" => rgb <= "100001";
                when "0100100101001" => rgb <= "100001";
                when "0100100101010" => rgb <= "100001";
                when "0100100101011" => rgb <= "100001";
                when "0100100101100" => rgb <= "100001";
                when "0100100101101" => rgb <= "100001";
                when "0100100110010" => rgb <= "100001";
                when "0100100110011" => rgb <= "100001";
                when "0100100110100" => rgb <= "100001";
                when "0100100110101" => rgb <= "100001";
                when "0100100110111" => rgb <= "100001";
                when "0100100111000" => rgb <= "100001";
                when "0100100111001" => rgb <= "010000";
                when "0100100111010" => rgb <= "010000";
                when "0100100111011" => rgb <= "100001";
                when "0100101000010" => rgb <= "100001";
                when "0100101000011" => rgb <= "100001";
                when "0100101000100" => rgb <= "100001";
                when "0100101000101" => rgb <= "100001";
                when "0100101000110" => rgb <= "010000";
                when "0100101000111" => rgb <= "100001";
                when "0100101001000" => rgb <= "100001";
                when "0100101001001" => rgb <= "100001";
                when "0100110001010" => rgb <= "100001";
                when "0100110001011" => rgb <= "100001";
                when "0100110001100" => rgb <= "010000";
                when "0100110001101" => rgb <= "100001";
                when "0100110010110" => rgb <= "100001";
                when "0100110010111" => rgb <= "100001";
                when "0100110011000" => rgb <= "100100";
                when "0100110011001" => rgb <= "100001";
                when "0100110011010" => rgb <= "010000";
                when "0100110011011" => rgb <= "010000";
                when "0100110011100" => rgb <= "010000";
                when "0100110011101" => rgb <= "100001";
                when "0100110011110" => rgb <= "100001";
                when "0100110011111" => rgb <= "100001";
                when "0100110100000" => rgb <= "100001";
                when "0100110100001" => rgb <= "100001";
                when "0100110100110" => rgb <= "010000";
                when "0100110100111" => rgb <= "100001";
                when "0100110101000" => rgb <= "100001";
                when "0100110101001" => rgb <= "100001";
                when "0100110101010" => rgb <= "100001";
                when "0100110101011" => rgb <= "100001";
                when "0100110101100" => rgb <= "100001";
                when "0100110101101" => rgb <= "100001";
                when "0100110110010" => rgb <= "100001";
                when "0100110110011" => rgb <= "100100";
                when "0100110110100" => rgb <= "100001";
                when "0100110110101" => rgb <= "100001";
                when "0100110111000" => rgb <= "100001";
                when "0100110111001" => rgb <= "100001";
                when "0100110111010" => rgb <= "100001";
                when "0100110111011" => rgb <= "100001";
                when "0100110111100" => rgb <= "100001";
                when "0100111000010" => rgb <= "100001";
                when "0100111000011" => rgb <= "100001";
                when "0100111000100" => rgb <= "100001";
                when "0100111000101" => rgb <= "100001";
                when "0100111000110" => rgb <= "100001";
                when "0100111000111" => rgb <= "100100";
                when "0100111001000" => rgb <= "100100";
                when "0100111001001" => rgb <= "100100";
                when "0101000001010" => rgb <= "100001";
                when "0101000001011" => rgb <= "100100";
                when "0101000001100" => rgb <= "100001";
                when "0101000001101" => rgb <= "010000";
                when "0101000011000" => rgb <= "100001";
                when "0101000011001" => rgb <= "100001";
                when "0101000011010" => rgb <= "100001";
                when "0101000011011" => rgb <= "100001";
                when "0101000011100" => rgb <= "100001";
                when "0101000011101" => rgb <= "100100";
                when "0101000011110" => rgb <= "100100";
                when "0101000011111" => rgb <= "100001";
                when "0101000100110" => rgb <= "100001";
                when "0101000100111" => rgb <= "001011";
                when "0101000101000" => rgb <= "100001";
                when "0101000101001" => rgb <= "010000";
                when "0101000101010" => rgb <= "100001";
                when "0101000101011" => rgb <= "100100";
                when "0101000101100" => rgb <= "100100";
                when "0101000101101" => rgb <= "100001";
                when "0101000110010" => rgb <= "100001";
                when "0101000110011" => rgb <= "100001";
                when "0101000110100" => rgb <= "100100";
                when "0101000110101" => rgb <= "100001";
                when "0101000111001" => rgb <= "100001";
                when "0101000111010" => rgb <= "100001";
                when "0101000111011" => rgb <= "100100";
                when "0101000111100" => rgb <= "100100";
                when "0101000111101" => rgb <= "100001";
                when "0101001000010" => rgb <= "100001";
                when "0101001000011" => rgb <= "100001";
                when "0101001000100" => rgb <= "100001";
                when "0101001000101" => rgb <= "100100";
                when "0101001000110" => rgb <= "100001";
                when "0101001000111" => rgb <= "100001";
                when "0101001001000" => rgb <= "100100";
                when "0101001001001" => rgb <= "100001";
                when "0101010001010" => rgb <= "010000";
                when "0101010001011" => rgb <= "100001";
                when "0101010001100" => rgb <= "100001";
                when "0101010001101" => rgb <= "100001";
                when "0101010011000" => rgb <= "100100";
                when "0101010011001" => rgb <= "100001";
                when "0101010011010" => rgb <= "100001";
                when "0101010011011" => rgb <= "100001";
                when "0101010011100" => rgb <= "010000";
                when "0101010011101" => rgb <= "100001";
                when "0101010011110" => rgb <= "100001";
                when "0101010011111" => rgb <= "100001";
                when "0101010100110" => rgb <= "100001";
                when "0101010100111" => rgb <= "001011";
                when "0101010101000" => rgb <= "100001";
                when "0101010101001" => rgb <= "100001";
                when "0101010101010" => rgb <= "010000";
                when "0101010101011" => rgb <= "010000";
                when "0101010101100" => rgb <= "010000";
                when "0101010101101" => rgb <= "100001";
                when "0101010110010" => rgb <= "100001";
                when "0101010110011" => rgb <= "100001";
                when "0101010110100" => rgb <= "100001";
                when "0101010110101" => rgb <= "100001";
                when "0101010111010" => rgb <= "010000";
                when "0101010111011" => rgb <= "010000";
                when "0101010111100" => rgb <= "100001";
                when "0101010111101" => rgb <= "100001";
                when "0101011000010" => rgb <= "010000";
                when "0101011000011" => rgb <= "100001";
                when "0101011000100" => rgb <= "100001";
                when "0101011000101" => rgb <= "100001";
                when "0101011000110" => rgb <= "100001";
                when "0101011000111" => rgb <= "100001";
                when "0101011001000" => rgb <= "100001";
                when "0101011001001" => rgb <= "100001";
                when "0110000010100" => rgb <= "111111";
                when "0110000010101" => rgb <= "111111";
                when "0110000010110" => rgb <= "111111";
                when "0110000011001" => rgb <= "111111";
                when "0110000011010" => rgb <= "111111";
                when "0110000011011" => rgb <= "111111";
                when "0110000011100" => rgb <= "111111";
                when "0110000011110" => rgb <= "111111";
                when "0110000011111" => rgb <= "111111";
                when "0110000100000" => rgb <= "111111";
                when "0110000100001" => rgb <= "111111";
                when "0110000100010" => rgb <= "111111";
                when "0110000100100" => rgb <= "111111";
                when "0110000100101" => rgb <= "111111";
                when "0110000100110" => rgb <= "111111";
                when "0110000101011" => rgb <= "111111";
                when "0110000101100" => rgb <= "111111";
                when "0110000101101" => rgb <= "111111";
                when "0110000101110" => rgb <= "111111";
                when "0110000110000" => rgb <= "111111";
                when "0110000110101" => rgb <= "111111";
                when "0110000110111" => rgb <= "111111";
                when "0110000111000" => rgb <= "111111";
                when "0110000111001" => rgb <= "111111";
                when "0110000111011" => rgb <= "111111";
                when "0110000111100" => rgb <= "111111";
                when "0110000111101" => rgb <= "111111";
                when "0110000111110" => rgb <= "111111";
                when "0110010010011" => rgb <= "111111";
                when "0110010010111" => rgb <= "111111";
                when "0110010011001" => rgb <= "111111";
                when "0110010011100" => rgb <= "111111";
                when "0110010011110" => rgb <= "111111";
                when "0110010100000" => rgb <= "111111";
                when "0110010100010" => rgb <= "111111";
                when "0110010100100" => rgb <= "111111";
                when "0110010101011" => rgb <= "111111";
                when "0110010101110" => rgb <= "111111";
                when "0110010110000" => rgb <= "111111";
                when "0110010110101" => rgb <= "111111";
                when "0110010110111" => rgb <= "111111";
                when "0110010111011" => rgb <= "111111";
                when "0110010111110" => rgb <= "111111";
                when "0110100010011" => rgb <= "111111";
                when "0110100011001" => rgb <= "111111";
                when "0110100011100" => rgb <= "111111";
                when "0110100011110" => rgb <= "111111";
                when "0110100100000" => rgb <= "111111";
                when "0110100100010" => rgb <= "111111";
                when "0110100100100" => rgb <= "111111";
                when "0110100101011" => rgb <= "111111";
                when "0110100101110" => rgb <= "111111";
                when "0110100110000" => rgb <= "111111";
                when "0110100110101" => rgb <= "111111";
                when "0110100110111" => rgb <= "111111";
                when "0110100111011" => rgb <= "111111";
                when "0110100111110" => rgb <= "111111";
                when "0110110010011" => rgb <= "111111";
                when "0110110011001" => rgb <= "111111";
                when "0110110011010" => rgb <= "111111";
                when "0110110011011" => rgb <= "111111";
                when "0110110011100" => rgb <= "111111";
                when "0110110011110" => rgb <= "111111";
                when "0110110100010" => rgb <= "111111";
                when "0110110100100" => rgb <= "111111";
                when "0110110100101" => rgb <= "111111";
                when "0110110100110" => rgb <= "111111";
                when "0110110101011" => rgb <= "111111";
                when "0110110101110" => rgb <= "111111";
                when "0110110110000" => rgb <= "111111";
                when "0110110110101" => rgb <= "111111";
                when "0110110110111" => rgb <= "111111";
                when "0110110111000" => rgb <= "111111";
                when "0110110111001" => rgb <= "111111";
                when "0110110111011" => rgb <= "111111";
                when "0110110111100" => rgb <= "111111";
                when "0110110111101" => rgb <= "111111";
                when "0110110111110" => rgb <= "111111";
                when "0111000010011" => rgb <= "111111";
                when "0111000010110" => rgb <= "111111";
                when "0111000010111" => rgb <= "111111";
                when "0111000011001" => rgb <= "111111";
                when "0111000011100" => rgb <= "111111";
                when "0111000011110" => rgb <= "111111";
                when "0111000100010" => rgb <= "111111";
                when "0111000100100" => rgb <= "111111";
                when "0111000101011" => rgb <= "111111";
                when "0111000101110" => rgb <= "111111";
                when "0111000110000" => rgb <= "111111";
                when "0111000110101" => rgb <= "111111";
                when "0111000110111" => rgb <= "111111";
                when "0111000111011" => rgb <= "111111";
                when "0111000111100" => rgb <= "111111";
                when "0111010010011" => rgb <= "111111";
                when "0111010010111" => rgb <= "111111";
                when "0111010011001" => rgb <= "111111";
                when "0111010011100" => rgb <= "111111";
                when "0111010011110" => rgb <= "111111";
                when "0111010100010" => rgb <= "111111";
                when "0111010100100" => rgb <= "111111";
                when "0111010101011" => rgb <= "111111";
                when "0111010101110" => rgb <= "111111";
                when "0111010110001" => rgb <= "111111";
                when "0111010110100" => rgb <= "111111";
                when "0111010110111" => rgb <= "111111";
                when "0111010111011" => rgb <= "111111";
                when "0111010111101" => rgb <= "111111";
                when "0111100010100" => rgb <= "111111";
                when "0111100010101" => rgb <= "111111";
                when "0111100010110" => rgb <= "111111";
                when "0111100010111" => rgb <= "111111";
                when "0111100011001" => rgb <= "111111";
                when "0111100011100" => rgb <= "111111";
                when "0111100011110" => rgb <= "111111";
                when "0111100100010" => rgb <= "111111";
                when "0111100100100" => rgb <= "111111";
                when "0111100100101" => rgb <= "111111";
                when "0111100100110" => rgb <= "111111";
                when "0111100101011" => rgb <= "111111";
                when "0111100101100" => rgb <= "111111";
                when "0111100101101" => rgb <= "111111";
                when "0111100101110" => rgb <= "111111";
                when "0111100110010" => rgb <= "111111";
                when "0111100110011" => rgb <= "111111";
                when "0111100110111" => rgb <= "111111";
                when "0111100111000" => rgb <= "111111";
                when "0111100111001" => rgb <= "111111";
                when "0111100111011" => rgb <= "111111";
                when "0111100111110" => rgb <= "111111";
                when "1000100011001" => rgb <= "001011";
                when "1000100011010" => rgb <= "001011";
                when "1000100011011" => rgb <= "001011";
                when "1000100011110" => rgb <= "001011";
                when "1000100100100" => rgb <= "001011";
                when "1000100100101" => rgb <= "001011";
                when "1000100101000" => rgb <= "001011";
                when "1000100101100" => rgb <= "001011";
                when "1000100101110" => rgb <= "001011";
                when "1000100101111" => rgb <= "001011";
                when "1000100110000" => rgb <= "001011";
                when "1000100110001" => rgb <= "001011";
                when "1000100110011" => rgb <= "001011";
                when "1000100110100" => rgb <= "001011";
                when "1000100110101" => rgb <= "001011";
                when "1000110011001" => rgb <= "001011";
                when "1000110011100" => rgb <= "001011";
                when "1000110011110" => rgb <= "001011";
                when "1000110100011" => rgb <= "001011";
                when "1000110100110" => rgb <= "001011";
                when "1000110101000" => rgb <= "001011";
                when "1000110101100" => rgb <= "001011";
                when "1000110101110" => rgb <= "001011";
                when "1000110110011" => rgb <= "001011";
                when "1000110110110" => rgb <= "001011";
                when "1001000011001" => rgb <= "001011";
                when "1001000011010" => rgb <= "001011";
                when "1001000011011" => rgb <= "001011";
                when "1001000011110" => rgb <= "001011";
                when "1001000100011" => rgb <= "001011";
                when "1001000100100" => rgb <= "001011";
                when "1001000100101" => rgb <= "001011";
                when "1001000100110" => rgb <= "001011";
                when "1001000101001" => rgb <= "001011";
                when "1001000101010" => rgb <= "001011";
                when "1001000101011" => rgb <= "001011";
                when "1001000101110" => rgb <= "001011";
                when "1001000101111" => rgb <= "001011";
                when "1001000110000" => rgb <= "001011";
                when "1001000110011" => rgb <= "001011";
                when "1001000110100" => rgb <= "001011";
                when "1001000110101" => rgb <= "001011";
                when "1001000111011" => rgb <= "010000";
                when "1001000111111" => rgb <= "111111";
                when "1001010011001" => rgb <= "001011";
                when "1001010011110" => rgb <= "001011";
                when "1001010100011" => rgb <= "001011";
                when "1001010100110" => rgb <= "001011";
                when "1001010101010" => rgb <= "001011";
                when "1001010101110" => rgb <= "001011";
                when "1001010110011" => rgb <= "001011";
                when "1001010110101" => rgb <= "001011";
                when "1001010111010" => rgb <= "111111";
                when "1001010111011" => rgb <= "010000";
                when "1001010111100" => rgb <= "010000";
                when "1001010111110" => rgb <= "111111";
                when "1001010111111" => rgb <= "111111";
                when "1001011000000" => rgb <= "111111";
                when "1001100001101" => rgb <= "111111";
                when "1001100001110" => rgb <= "111111";
                when "1001100001111" => rgb <= "111111";
                when "1001100010000" => rgb <= "111111";
                when "1001100010001" => rgb <= "111111";
                when "1001100010010" => rgb <= "111111";
                when "1001100010011" => rgb <= "111111";
                when "1001100010100" => rgb <= "111111";
                when "1001100010101" => rgb <= "111111";
                when "1001100010110" => rgb <= "111111";
                when "1001100011001" => rgb <= "001011";
                when "1001100011110" => rgb <= "001011";
                when "1001100011111" => rgb <= "001011";
                when "1001100100000" => rgb <= "001011";
                when "1001100100001" => rgb <= "001011";
                when "1001100100011" => rgb <= "001011";
                when "1001100100110" => rgb <= "001011";
                when "1001100101010" => rgb <= "001011";
                when "1001100101110" => rgb <= "001011";
                when "1001100101111" => rgb <= "001011";
                when "1001100110000" => rgb <= "001011";
                when "1001100110001" => rgb <= "001011";
                when "1001100110011" => rgb <= "001011";
                when "1001100110110" => rgb <= "001011";
                when "1001100111010" => rgb <= "111111";
                when "1001100111011" => rgb <= "010000";
                when "1001100111100" => rgb <= "111111";
                when "1001100111101" => rgb <= "111111";
                when "1001100111110" => rgb <= "111111";
                when "1001100111111" => rgb <= "111111";
                when "1001101000000" => rgb <= "111111";
                when "1001110001101" => rgb <= "111111";
                when "1001110001110" => rgb <= "111111";
                when "1001110001111" => rgb <= "111111";
                when "1001110010000" => rgb <= "111111";
                when "1001110010001" => rgb <= "111111";
                when "1001110010010" => rgb <= "111111";
                when "1001110010011" => rgb <= "111111";
                when "1001110010100" => rgb <= "111111";
                when "1001110010101" => rgb <= "111111";
                when "1001110010110" => rgb <= "111111";
                when "1001110111011" => rgb <= "111111";
                when "1001110111100" => rgb <= "111111";
                when "1001110111101" => rgb <= "010000";
                when "1001110111110" => rgb <= "111111";
                when "1001110111111" => rgb <= "111111";
                when "1010000000111" => rgb <= "111111";
                when "1010000001000" => rgb <= "111111";
                when "1010000001001" => rgb <= "111111";
                when "1010000001010" => rgb <= "111111";
                when "1010000001011" => rgb <= "111111";
                when "1010000001100" => rgb <= "111111";
                when "1010000001101" => rgb <= "111111";
                when "1010000001110" => rgb <= "111111";
                when "1010000001111" => rgb <= "111111";
                when "1010000010000" => rgb <= "111111";
                when "1010000010001" => rgb <= "111111";
                when "1010000010010" => rgb <= "111111";
                when "1010000010011" => rgb <= "111111";
                when "1010000010100" => rgb <= "111111";
                when "1010000010101" => rgb <= "111111";
                when "1010000010110" => rgb <= "111111";
                when "1010000010111" => rgb <= "111111";
                when "1010000011000" => rgb <= "111111";
                when "1010000111100" => rgb <= "010000";
                when "1010000111101" => rgb <= "010000";
                when "1010000111110" => rgb <= "111111";
                when "1010001000011" => rgb <= "111111";
                when "1010001000100" => rgb <= "111111";
                when "1010001000101" => rgb <= "111111";
                when "1010001000110" => rgb <= "111111";
                when "1010001000111" => rgb <= "111111";
                when "1010001001000" => rgb <= "111111";
                when "1010010000111" => rgb <= "111111";
                when "1010010001000" => rgb <= "111111";
                when "1010010001001" => rgb <= "111111";
                when "1010010001010" => rgb <= "111111";
                when "1010010001011" => rgb <= "111111";
                when "1010010001100" => rgb <= "111111";
                when "1010010001101" => rgb <= "111111";
                when "1010010001110" => rgb <= "111111";
                when "1010010001111" => rgb <= "111111";
                when "1010010010000" => rgb <= "111111";
                when "1010010010001" => rgb <= "111111";
                when "1010010010010" => rgb <= "111111";
                when "1010010010011" => rgb <= "111111";
                when "1010010010100" => rgb <= "111111";
                when "1010010010101" => rgb <= "111111";
                when "1010010010110" => rgb <= "111111";
                when "1010010010111" => rgb <= "111111";
                when "1010010011000" => rgb <= "111111";
                when "1010010101000" => rgb <= "001011";
                when "1010010111100" => rgb <= "111111";
                when "1010010111101" => rgb <= "010000";
                when "1010010111110" => rgb <= "111111";
                when "1010011000010" => rgb <= "111111";
                when "1010011000011" => rgb <= "111111";
                when "1010011000100" => rgb <= "111111";
                when "1010011000101" => rgb <= "111111";
                when "1010011000110" => rgb <= "111111";
                when "1010011000111" => rgb <= "111111";
                when "1010011001000" => rgb <= "111111";
                when "1010100000101" => rgb <= "111111";
                when "1010100000110" => rgb <= "111111";
                when "1010100000111" => rgb <= "111111";
                when "1010100001000" => rgb <= "111111";
                when "1010100001001" => rgb <= "111111";
                when "1010100001010" => rgb <= "111111";
                when "1010100001011" => rgb <= "111111";
                when "1010100001100" => rgb <= "111111";
                when "1010100001101" => rgb <= "111111";
                when "1010100001110" => rgb <= "111111";
                when "1010100001111" => rgb <= "111111";
                when "1010100010000" => rgb <= "111111";
                when "1010100010001" => rgb <= "111111";
                when "1010100010010" => rgb <= "111111";
                when "1010100010011" => rgb <= "111111";
                when "1010100010100" => rgb <= "111111";
                when "1010100010101" => rgb <= "111111";
                when "1010100010110" => rgb <= "111111";
                when "1010100010111" => rgb <= "111111";
                when "1010100011000" => rgb <= "111111";
                when "1010100100111" => rgb <= "001011";
                when "1010100101000" => rgb <= "001011";
                when "1010100111100" => rgb <= "111111";
                when "1010100111101" => rgb <= "111111";
                when "1010100111110" => rgb <= "010000";
                when "1010101000001" => rgb <= "111111";
                when "1010101000010" => rgb <= "111111";
                when "1010101000011" => rgb <= "111111";
                when "1010101000100" => rgb <= "111111";
                when "1010101000101" => rgb <= "111111";
                when "1010101000110" => rgb <= "111111";
                when "1010101000111" => rgb <= "111111";
                when "1010101001000" => rgb <= "111111";
                when "1010101001001" => rgb <= "111111";
                when "1010101001010" => rgb <= "111111";
                when "1010110000101" => rgb <= "111111";
                when "1010110000110" => rgb <= "111111";
                when "1010110000111" => rgb <= "111111";
                when "1010110001000" => rgb <= "111111";
                when "1010110001001" => rgb <= "111111";
                when "1010110001010" => rgb <= "111111";
                when "1010110001011" => rgb <= "111111";
                when "1010110001100" => rgb <= "111111";
                when "1010110001101" => rgb <= "111111";
                when "1010110001110" => rgb <= "111111";
                when "1010110001111" => rgb <= "111111";
                when "1010110010000" => rgb <= "111111";
                when "1010110010001" => rgb <= "111111";
                when "1010110010010" => rgb <= "111111";
                when "1010110010011" => rgb <= "111111";
                when "1010110010100" => rgb <= "111111";
                when "1010110010101" => rgb <= "111111";
                when "1010110010110" => rgb <= "111111";
                when "1010110010111" => rgb <= "111111";
                when "1010110011000" => rgb <= "111111";
                when "1010110101000" => rgb <= "001011";
                when "1010110111100" => rgb <= "111111";
                when "1010110111101" => rgb <= "010000";
                when "1010110111110" => rgb <= "010000";
                when "1010111000000" => rgb <= "111111";
                when "1010111000001" => rgb <= "111111";
                when "1010111000010" => rgb <= "111111";
                when "1010111000011" => rgb <= "111111";
                when "1010111000100" => rgb <= "111111";
                when "1010111000101" => rgb <= "111111";
                when "1010111000110" => rgb <= "111111";
                when "1010111000111" => rgb <= "111111";
                when "1010111001000" => rgb <= "111111";
                when "1010111001001" => rgb <= "111111";
                when "1010111001010" => rgb <= "111111";
                when "1011000000011" => rgb <= "111111";
                when "1011000000100" => rgb <= "111111";
                when "1011000000101" => rgb <= "111111";
                when "1011000000110" => rgb <= "111111";
                when "1011000000111" => rgb <= "111111";
                when "1011000001000" => rgb <= "111111";
                when "1011000001001" => rgb <= "111111";
                when "1011000001010" => rgb <= "111111";
                when "1011000001011" => rgb <= "111111";
                when "1011000001100" => rgb <= "111111";
                when "1011000001101" => rgb <= "111111";
                when "1011000001110" => rgb <= "111111";
                when "1011000001111" => rgb <= "111111";
                when "1011000010000" => rgb <= "111111";
                when "1011000010001" => rgb <= "111111";
                when "1011000010010" => rgb <= "111111";
                when "1011000010101" => rgb <= "111111";
                when "1011000010110" => rgb <= "111111";
                when "1011000010111" => rgb <= "111111";
                when "1011000011000" => rgb <= "111111";
                when "1011000101000" => rgb <= "001011";
                when "1011000111100" => rgb <= "111111";
                when "1011000111101" => rgb <= "010000";
                when "1011000111110" => rgb <= "101010";
                when "1011000111111" => rgb <= "010000";
                when "1011001000000" => rgb <= "111111";
                when "1011001000001" => rgb <= "111111";
                when "1011001000010" => rgb <= "111111";
                when "1011001000011" => rgb <= "111111";
                when "1011001000100" => rgb <= "111111";
                when "1011001000101" => rgb <= "111111";
                when "1011001000110" => rgb <= "111111";
                when "1011001000111" => rgb <= "111111";
                when "1011001001000" => rgb <= "111111";
                when "1011001001001" => rgb <= "111111";
                when "1011001001010" => rgb <= "111111";
                when "1011001001011" => rgb <= "111111";
                when "1011001001100" => rgb <= "111111";
                when "1011010000011" => rgb <= "111111";
                when "1011010000100" => rgb <= "111111";
                when "1011010000101" => rgb <= "111111";
                when "1011010000110" => rgb <= "111111";
                when "1011010000111" => rgb <= "111111";
                when "1011010001000" => rgb <= "111111";
                when "1011010001001" => rgb <= "111111";
                when "1011010001010" => rgb <= "111111";
                when "1011010001011" => rgb <= "111111";
                when "1011010001100" => rgb <= "111111";
                when "1011010001101" => rgb <= "111111";
                when "1011010001110" => rgb <= "111111";
                when "1011010001111" => rgb <= "111111";
                when "1011010010000" => rgb <= "111111";
                when "1011010010001" => rgb <= "111111";
                when "1011010010010" => rgb <= "111111";
                when "1011010010101" => rgb <= "111111";
                when "1011010010110" => rgb <= "111111";
                when "1011010010111" => rgb <= "111111";
                when "1011010011000" => rgb <= "111111";
                when "1011010100111" => rgb <= "001011";
                when "1011010101000" => rgb <= "001011";
                when "1011010101001" => rgb <= "001011";
                when "1011010111100" => rgb <= "111111";
                when "1011010111101" => rgb <= "101010";
                when "1011010111110" => rgb <= "010000";
                when "1011010111111" => rgb <= "111111";
                when "1011011000000" => rgb <= "010000";
                when "1011011000001" => rgb <= "111111";
                when "1011011000010" => rgb <= "111111";
                when "1011011000011" => rgb <= "111111";
                when "1011011000100" => rgb <= "111111";
                when "1011011000101" => rgb <= "111111";
                when "1011011000110" => rgb <= "111111";
                when "1011011000111" => rgb <= "111111";
                when "1011011001000" => rgb <= "111111";
                when "1011011001001" => rgb <= "111111";
                when "1011011001010" => rgb <= "111111";
                when "1011011001011" => rgb <= "111111";
                when "1011011001100" => rgb <= "111111";
                when "1011100000001" => rgb <= "111111";
                when "1011100000010" => rgb <= "111111";
                when "1011100000011" => rgb <= "111111";
                when "1011100000100" => rgb <= "111111";
                when "1011100000101" => rgb <= "111111";
                when "1011100000110" => rgb <= "111111";
                when "1011100000111" => rgb <= "111111";
                when "1011100001000" => rgb <= "111111";
                when "1011100001001" => rgb <= "111111";
                when "1011100001010" => rgb <= "111111";
                when "1011100001011" => rgb <= "111111";
                when "1011100001100" => rgb <= "111111";
                when "1011100001101" => rgb <= "111111";
                when "1011100001110" => rgb <= "111111";
                when "1011100001111" => rgb <= "111111";
                when "1011100010000" => rgb <= "111111";
                when "1011100010001" => rgb <= "111111";
                when "1011100010010" => rgb <= "111111";
                when "1011100010011" => rgb <= "111111";
                when "1011100010100" => rgb <= "111111";
                when "1011100010101" => rgb <= "111111";
                when "1011100010110" => rgb <= "111111";
                when "1011100010111" => rgb <= "111111";
                when "1011100011000" => rgb <= "111111";
                when "1011100111100" => rgb <= "101010";
                when "1011100111101" => rgb <= "010000";
                when "1011100111110" => rgb <= "010000";
                when "1011100111111" => rgb <= "111111";
                when "1011101000000" => rgb <= "111111";
                when "1011101000001" => rgb <= "111111";
                when "1011101000010" => rgb <= "111111";
                when "1011101000011" => rgb <= "111111";
                when "1011101000100" => rgb <= "111111";
                when "1011101000101" => rgb <= "111111";
                when "1011101000110" => rgb <= "111111";
                when "1011101000111" => rgb <= "111111";
                when "1011101001000" => rgb <= "111111";
                when "1011101001001" => rgb <= "111111";
                when "1011101001010" => rgb <= "111111";
                when "1011101001011" => rgb <= "111111";
                when "1011101001100" => rgb <= "111111";
                when "1011101001101" => rgb <= "111111";
                when "1011101001110" => rgb <= "111111";
                when "1011110000001" => rgb <= "111111";
                when "1011110000010" => rgb <= "111111";
                when "1011110000011" => rgb <= "111111";
                when "1011110000100" => rgb <= "111111";
                when "1011110000101" => rgb <= "111111";
                when "1011110000110" => rgb <= "111111";
                when "1011110000111" => rgb <= "111111";
                when "1011110001000" => rgb <= "111111";
                when "1011110001001" => rgb <= "111111";
                when "1011110001010" => rgb <= "111111";
                when "1011110001011" => rgb <= "111111";
                when "1011110001100" => rgb <= "111111";
                when "1011110001101" => rgb <= "111111";
                when "1011110001110" => rgb <= "111111";
                when "1011110001111" => rgb <= "111111";
                when "1011110010000" => rgb <= "111111";
                when "1011110010001" => rgb <= "111111";
                when "1011110010010" => rgb <= "111111";
                when "1011110010011" => rgb <= "111111";
                when "1011110010100" => rgb <= "111111";
                when "1011110010101" => rgb <= "111111";
                when "1011110010110" => rgb <= "111111";
                when "1011110010111" => rgb <= "111111";
                when "1011110011000" => rgb <= "111111";
                when "1011110111100" => rgb <= "010000";
                when "1011110111101" => rgb <= "111111";
                when "1011110111110" => rgb <= "010000";
                when "1011110111111" => rgb <= "111111";
                when "1011111000000" => rgb <= "111111";
                when "1011111000001" => rgb <= "111111";
                when "1011111000010" => rgb <= "111111";
                when "1011111000011" => rgb <= "111111";
                when "1011111000100" => rgb <= "111111";
                when "1011111000101" => rgb <= "111111";
                when "1011111000110" => rgb <= "111111";
                when "1011111000111" => rgb <= "111111";
                when "1011111001000" => rgb <= "111111";
                when "1011111001001" => rgb <= "111111";
                when "1011111001010" => rgb <= "111111";
                when "1011111001011" => rgb <= "111111";
                when "1011111001100" => rgb <= "111111";
                when "1011111001101" => rgb <= "111111";
                when "1011111001110" => rgb <= "111111";
                when "1100000000011" => rgb <= "111111";
                when "1100000000100" => rgb <= "111111";
                when "1100000000101" => rgb <= "111111";
                when "1100000000110" => rgb <= "111111";
                when "1100000000111" => rgb <= "111111";
                when "1100000001000" => rgb <= "111111";
                when "1100000001001" => rgb <= "111111";
                when "1100000001010" => rgb <= "111111";
                when "1100000001011" => rgb <= "111111";
                when "1100000001100" => rgb <= "111111";
                when "1100000001101" => rgb <= "111111";
                when "1100000001110" => rgb <= "111111";
                when "1100000001111" => rgb <= "111111";
                when "1100000010000" => rgb <= "111111";
                when "1100000010001" => rgb <= "111111";
                when "1100000010010" => rgb <= "111111";
                when "1100000010011" => rgb <= "111111";
                when "1100000010100" => rgb <= "111111";
                when "1100000010101" => rgb <= "111111";
                when "1100000010110" => rgb <= "111111";
                when "1100000010111" => rgb <= "111111";
                when "1100000011000" => rgb <= "111111";
                when "1100000011111" => rgb <= "001011";
                when "1100000100011" => rgb <= "001011";
                when "1100000100101" => rgb <= "001011";
                when "1100000100110" => rgb <= "001011";
                when "1100000100111" => rgb <= "001011";
                when "1100000101001" => rgb <= "001011";
                when "1100000101100" => rgb <= "001011";
                when "1100000101111" => rgb <= "001011";
                when "1100000110000" => rgb <= "001011";
                when "1100000110001" => rgb <= "001011";
                when "1100000111011" => rgb <= "010000";
                when "1100000111100" => rgb <= "010000";
                when "1100000111101" => rgb <= "111111";
                when "1100000111110" => rgb <= "111111";
                when "1100000111111" => rgb <= "111111";
                when "1100001000000" => rgb <= "111111";
                when "1100001000001" => rgb <= "111111";
                when "1100001000010" => rgb <= "111111";
                when "1100001000011" => rgb <= "111111";
                when "1100001000100" => rgb <= "111111";
                when "1100001000101" => rgb <= "111111";
                when "1100001000110" => rgb <= "111111";
                when "1100001000111" => rgb <= "111111";
                when "1100001001000" => rgb <= "111111";
                when "1100001001001" => rgb <= "111111";
                when "1100001001010" => rgb <= "111111";
                when "1100001001011" => rgb <= "111111";
                when "1100001001100" => rgb <= "111111";
                when "1100010000011" => rgb <= "111111";
                when "1100010000100" => rgb <= "111111";
                when "1100010000101" => rgb <= "111111";
                when "1100010000110" => rgb <= "111111";
                when "1100010000111" => rgb <= "111111";
                when "1100010001000" => rgb <= "111111";
                when "1100010001001" => rgb <= "111111";
                when "1100010001010" => rgb <= "111111";
                when "1100010001011" => rgb <= "111111";
                when "1100010001100" => rgb <= "111111";
                when "1100010001101" => rgb <= "111111";
                when "1100010001110" => rgb <= "111111";
                when "1100010001111" => rgb <= "111111";
                when "1100010010000" => rgb <= "111111";
                when "1100010010001" => rgb <= "111111";
                when "1100010010010" => rgb <= "111111";
                when "1100010010011" => rgb <= "111111";
                when "1100010010100" => rgb <= "111111";
                when "1100010010101" => rgb <= "111111";
                when "1100010010110" => rgb <= "111111";
                when "1100010010111" => rgb <= "111111";
                when "1100010011000" => rgb <= "111111";
                when "1100010011111" => rgb <= "001011";
                when "1100010100011" => rgb <= "001011";
                when "1100010100110" => rgb <= "001011";
                when "1100010101001" => rgb <= "001011";
                when "1100010101010" => rgb <= "001011";
                when "1100010101100" => rgb <= "001011";
                when "1100010101110" => rgb <= "001011";
                when "1100010111010" => rgb <= "111111";
                when "1100010111011" => rgb <= "010000";
                when "1100010111100" => rgb <= "111111";
                when "1100010111101" => rgb <= "111111";
                when "1100010111110" => rgb <= "111111";
                when "1100010111111" => rgb <= "111111";
                when "1100011000000" => rgb <= "111111";
                when "1100011000001" => rgb <= "111111";
                when "1100011000010" => rgb <= "111111";
                when "1100011000011" => rgb <= "111111";
                when "1100011000100" => rgb <= "111111";
                when "1100011000101" => rgb <= "111111";
                when "1100011000110" => rgb <= "111111";
                when "1100011000111" => rgb <= "111111";
                when "1100011001000" => rgb <= "111111";
                when "1100011001001" => rgb <= "111111";
                when "1100011001010" => rgb <= "111111";
                when "1100011001011" => rgb <= "111111";
                when "1100011001100" => rgb <= "111111";
                when "1100100000011" => rgb <= "111111";
                when "1100100000100" => rgb <= "111111";
                when "1100100000101" => rgb <= "111111";
                when "1100100000110" => rgb <= "111111";
                when "1100100000111" => rgb <= "111111";
                when "1100100001000" => rgb <= "111111";
                when "1100100001001" => rgb <= "111111";
                when "1100100001010" => rgb <= "111111";
                when "1100100001011" => rgb <= "111111";
                when "1100100001100" => rgb <= "111111";
                when "1100100001101" => rgb <= "111111";
                when "1100100001110" => rgb <= "111111";
                when "1100100001111" => rgb <= "111111";
                when "1100100010000" => rgb <= "111111";
                when "1100100010001" => rgb <= "111111";
                when "1100100010010" => rgb <= "111111";
                when "1100100010011" => rgb <= "111111";
                when "1100100010100" => rgb <= "111111";
                when "1100100010101" => rgb <= "111111";
                when "1100100010110" => rgb <= "111111";
                when "1100100010111" => rgb <= "111111";
                when "1100100011000" => rgb <= "111111";
                when "1100100011111" => rgb <= "001011";
                when "1100100100001" => rgb <= "001011";
                when "1100100100011" => rgb <= "001011";
                when "1100100100110" => rgb <= "001011";
                when "1100100101001" => rgb <= "001011";
                when "1100100101011" => rgb <= "001011";
                when "1100100101100" => rgb <= "001011";
                when "1100100101111" => rgb <= "001011";
                when "1100100110000" => rgb <= "001011";
                when "1100100111001" => rgb <= "111111";
                when "1100100111010" => rgb <= "111111";
                when "1100100111011" => rgb <= "010000";
                when "1100100111100" => rgb <= "111111";
                when "1100100111101" => rgb <= "111111";
                when "1100100111110" => rgb <= "111111";
                when "1100100111111" => rgb <= "111111";
                when "1100101000000" => rgb <= "111111";
                when "1100101000001" => rgb <= "111111";
                when "1100101000010" => rgb <= "111111";
                when "1100101000011" => rgb <= "111111";
                when "1100101000100" => rgb <= "111111";
                when "1100101000101" => rgb <= "111111";
                when "1100101000110" => rgb <= "111111";
                when "1100101000111" => rgb <= "111111";
                when "1100101001000" => rgb <= "111111";
                when "1100101001001" => rgb <= "111111";
                when "1100101001010" => rgb <= "111111";
                when "1100101001011" => rgb <= "111111";
                when "1100101001100" => rgb <= "111111";
                when "1100110000011" => rgb <= "111111";
                when "1100110000100" => rgb <= "111111";
                when "1100110000101" => rgb <= "111111";
                when "1100110000110" => rgb <= "111111";
                when "1100110000111" => rgb <= "111111";
                when "1100110001000" => rgb <= "111111";
                when "1100110001001" => rgb <= "111111";
                when "1100110001010" => rgb <= "111111";
                when "1100110001011" => rgb <= "111111";
                when "1100110001100" => rgb <= "111111";
                when "1100110001101" => rgb <= "111111";
                when "1100110001110" => rgb <= "111111";
                when "1100110001111" => rgb <= "111111";
                when "1100110010000" => rgb <= "111111";
                when "1100110010001" => rgb <= "111111";
                when "1100110010010" => rgb <= "111111";
                when "1100110010011" => rgb <= "111111";
                when "1100110010100" => rgb <= "111111";
                when "1100110010101" => rgb <= "111111";
                when "1100110010110" => rgb <= "111111";
                when "1100110010111" => rgb <= "111111";
                when "1100110011000" => rgb <= "111111";
                when "1100110011111" => rgb <= "001011";
                when "1100110100000" => rgb <= "001011";
                when "1100110100010" => rgb <= "001011";
                when "1100110100011" => rgb <= "001011";
                when "1100110100110" => rgb <= "001011";
                when "1100110101001" => rgb <= "001011";
                when "1100110101100" => rgb <= "001011";
                when "1100110110001" => rgb <= "001011";
                when "1100110111000" => rgb <= "111111";
                when "1100110111001" => rgb <= "111111";
                when "1100110111010" => rgb <= "111111";
                when "1100110111011" => rgb <= "111111";
                when "1100110111100" => rgb <= "111111";
                when "1100110111101" => rgb <= "111111";
                when "1100110111110" => rgb <= "111111";
                when "1100110111111" => rgb <= "111111";
                when "1100111000000" => rgb <= "111111";
                when "1100111000001" => rgb <= "111111";
                when "1100111000010" => rgb <= "111111";
                when "1100111000011" => rgb <= "111111";
                when "1100111000100" => rgb <= "111111";
                when "1100111000101" => rgb <= "111111";
                when "1100111000110" => rgb <= "111111";
                when "1100111000111" => rgb <= "111111";
                when "1100111001000" => rgb <= "111111";
                when "1100111001001" => rgb <= "111111";
                when "1100111001010" => rgb <= "111111";
                when "1100111001011" => rgb <= "111111";
                when "1100111001100" => rgb <= "111111";
                when "1101000000011" => rgb <= "111111";
                when "1101000000100" => rgb <= "111111";
                when "1101000000101" => rgb <= "111111";
                when "1101000000110" => rgb <= "111111";
                when "1101000000111" => rgb <= "111111";
                when "1101000001000" => rgb <= "111111";
                when "1101000001101" => rgb <= "111111";
                when "1101000001110" => rgb <= "111111";
                when "1101000001111" => rgb <= "111111";
                when "1101000010000" => rgb <= "111111";
                when "1101000010001" => rgb <= "111111";
                when "1101000010010" => rgb <= "111111";
                when "1101000010101" => rgb <= "111111";
                when "1101000010110" => rgb <= "111111";
                when "1101000010111" => rgb <= "111111";
                when "1101000011000" => rgb <= "111111";
                when "1101000011001" => rgb <= "111111";
                when "1101000011010" => rgb <= "111111";
                when "1101000011111" => rgb <= "001011";
                when "1101000100011" => rgb <= "001011";
                when "1101000100101" => rgb <= "001011";
                when "1101000100110" => rgb <= "001011";
                when "1101000100111" => rgb <= "001011";
                when "1101000101001" => rgb <= "001011";
                when "1101000101100" => rgb <= "001011";
                when "1101000101110" => rgb <= "001011";
                when "1101000101111" => rgb <= "001011";
                when "1101000110000" => rgb <= "001011";
                when "1101000111101" => rgb <= "111111";
                when "1101000111110" => rgb <= "111111";
                when "1101000111111" => rgb <= "111111";
                when "1101001000000" => rgb <= "111111";
                when "1101001000001" => rgb <= "111111";
                when "1101001000010" => rgb <= "111111";
                when "1101001000111" => rgb <= "111111";
                when "1101001001000" => rgb <= "111111";
                when "1101001001001" => rgb <= "111111";
                when "1101001001010" => rgb <= "111111";
                when "1101001001011" => rgb <= "111111";
                when "1101001001100" => rgb <= "111111";
                when "1101010000011" => rgb <= "111111";
                when "1101010000100" => rgb <= "111111";
                when "1101010000101" => rgb <= "111111";
                when "1101010000110" => rgb <= "111111";
                when "1101010000111" => rgb <= "111111";
                when "1101010001000" => rgb <= "111111";
                when "1101010001101" => rgb <= "111111";
                when "1101010001110" => rgb <= "111111";
                when "1101010001111" => rgb <= "111111";
                when "1101010010000" => rgb <= "111111";
                when "1101010010001" => rgb <= "111111";
                when "1101010010010" => rgb <= "111111";
                when "1101010010101" => rgb <= "111111";
                when "1101010010110" => rgb <= "111111";
                when "1101010010111" => rgb <= "111111";
                when "1101010011000" => rgb <= "111111";
                when "1101010011001" => rgb <= "111111";
                when "1101010011010" => rgb <= "111111";
                when "1101010111101" => rgb <= "111111";
                when "1101010111110" => rgb <= "111111";
                when "1101010111111" => rgb <= "111111";
                when "1101011000000" => rgb <= "111111";
                when "1101011000001" => rgb <= "111111";
                when "1101011000010" => rgb <= "111111";
                when "1101011000111" => rgb <= "111111";
                when "1101011001000" => rgb <= "111111";
                when "1101011001001" => rgb <= "111111";
                when "1101011001010" => rgb <= "111111";
                when "1101011001011" => rgb <= "111111";
                when "1101011001100" => rgb <= "111111";
                when "1101100000011" => rgb <= "111111";
                when "1101100000100" => rgb <= "111111";
                when "1101100000101" => rgb <= "111111";
                when "1101100000110" => rgb <= "111111";
                when "1101100000111" => rgb <= "111111";
                when "1101100001000" => rgb <= "111111";
                when "1101100001101" => rgb <= "111111";
                when "1101100001110" => rgb <= "111111";
                when "1101100001111" => rgb <= "111111";
                when "1101100010000" => rgb <= "111111";
                when "1101100010001" => rgb <= "111111";
                when "1101100010010" => rgb <= "111111";
                when "1101100011001" => rgb <= "111111";
                when "1101100011010" => rgb <= "111111";
                when "1101100011011" => rgb <= "111111";
                when "1101100011100" => rgb <= "111111";
                when "1101100111101" => rgb <= "111111";
                when "1101100111110" => rgb <= "111111";
                when "1101100111111" => rgb <= "111111";
                when "1101101000000" => rgb <= "111111";
                when "1101101000001" => rgb <= "111111";
                when "1101101000010" => rgb <= "111111";
                when "1101101000111" => rgb <= "111111";
                when "1101101001000" => rgb <= "111111";
                when "1101101001001" => rgb <= "111111";
                when "1101101001010" => rgb <= "111111";
                when "1101101001011" => rgb <= "111111";
                when "1101101001100" => rgb <= "111111";
                when "1101110000011" => rgb <= "111111";
                when "1101110000100" => rgb <= "111111";
                when "1101110000101" => rgb <= "111111";
                when "1101110000110" => rgb <= "111111";
                when "1101110000111" => rgb <= "111111";
                when "1101110001000" => rgb <= "111111";
                when "1101110001101" => rgb <= "111111";
                when "1101110001110" => rgb <= "111111";
                when "1101110001111" => rgb <= "111111";
                when "1101110010000" => rgb <= "111111";
                when "1101110010001" => rgb <= "111111";
                when "1101110010010" => rgb <= "111111";
                when "1101110011001" => rgb <= "111111";
                when "1101110011010" => rgb <= "111111";
                when "1101110011011" => rgb <= "111111";
                when "1101110011100" => rgb <= "111111";
                when "1101110111101" => rgb <= "111111";
                when "1101110111110" => rgb <= "111111";
                when "1101110111111" => rgb <= "111111";
                when "1101111000000" => rgb <= "111111";
                when "1101111000001" => rgb <= "111111";
                when "1101111000010" => rgb <= "111111";
                when "1101111000111" => rgb <= "111111";
                when "1101111001000" => rgb <= "111111";
                when "1101111001001" => rgb <= "111111";
                when "1101111001010" => rgb <= "111111";
                when "1101111001011" => rgb <= "111111";
                when "1101111001100" => rgb <= "111111";
                when "1110000000011" => rgb <= "111111";
                when "1110000000100" => rgb <= "111111";
                when "1110000000101" => rgb <= "111111";
                when "1110000000110" => rgb <= "111111";
                when "1110000000111" => rgb <= "111111";
                when "1110000001000" => rgb <= "111111";
                when "1110000001101" => rgb <= "111111";
                when "1110000001110" => rgb <= "111111";
                when "1110000001111" => rgb <= "111111";
                when "1110000010000" => rgb <= "111111";
                when "1110000010001" => rgb <= "111111";
                when "1110000010010" => rgb <= "111111";
                when "1110000111101" => rgb <= "111111";
                when "1110000111110" => rgb <= "111111";
                when "1110000111111" => rgb <= "111111";
                when "1110001000000" => rgb <= "111111";
                when "1110001000001" => rgb <= "111111";
                when "1110001000010" => rgb <= "111111";
                when "1110001000111" => rgb <= "111111";
                when "1110001001000" => rgb <= "111111";
                when "1110001001001" => rgb <= "111111";
                when "1110001001010" => rgb <= "111111";
                when "1110001001011" => rgb <= "111111";
                when "1110001001100" => rgb <= "111111";
                when "1110010000011" => rgb <= "111111";
                when "1110010000100" => rgb <= "111111";
                when "1110010000101" => rgb <= "111111";
                when "1110010000110" => rgb <= "111111";
                when "1110010000111" => rgb <= "111111";
                when "1110010001000" => rgb <= "111111";
                when "1110010001101" => rgb <= "111111";
                when "1110010001110" => rgb <= "111111";
                when "1110010001111" => rgb <= "111111";
                when "1110010010000" => rgb <= "111111";
                when "1110010010001" => rgb <= "111111";
                when "1110010010010" => rgb <= "111111";
                when "1110010111101" => rgb <= "111111";
                when "1110010111110" => rgb <= "111111";
                when "1110010111111" => rgb <= "111111";
                when "1110011000000" => rgb <= "111111";
                when "1110011000001" => rgb <= "111111";
                when "1110011000010" => rgb <= "111111";
                when "1110011000111" => rgb <= "111111";
                when "1110011001000" => rgb <= "111111";
                when "1110011001001" => rgb <= "111111";
                when "1110011001010" => rgb <= "111111";
                when "1110011001011" => rgb <= "111111";
                when "1110011001100" => rgb <= "111111";
                when others => rgb <= "000000";
			end case;
		end if;
	end process;
	location <= std_logic_vector(col_idx) & std_logic_vector(row_idx);
end;