library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity start_rom is
  port(
	  clk : in std_logic;
	  row_idx: in unsigned(6 downto 0);
	  col_idx : in unsigned(5 downto 0); 
	  rgb : out std_logic_vector(5 downto 0)
	  );
end start_rom;

architecture synth of start_rom is

signal location : std_logic_vector(12 downto 0);
begin
	process (clk) begin
		if rising_edge(clk) then
			case location is
				when "0010000000110" => rgb <= "100001";
				when "0010000000111" => rgb <= "100100";
				when "0010000001000" => rgb <= "100100";
				when "0010000001001" => rgb <= "100100";
				when "0010000001010" => rgb <= "100100";
				when "0010000001011" => rgb <= "100001";
				when "0010000001100" => rgb <= "100001";
				when "0010000001101" => rgb <= "100001";
				when "0010000001110" => rgb <= "100001";
				when "0010000001111" => rgb <= "010000";
				when "0010000010000" => rgb <= "100001";
				when "0010000010001" => rgb <= "100001";
				when "0010000010110" => rgb <= "100001";
				when "0010000010111" => rgb <= "100001";
				when "0010000011000" => rgb <= "100001";
				when "0010000011001" => rgb <= "100100";
				when "0010000011110" => rgb <= "100001";
				when "0010000011111" => rgb <= "100001";
				when "0010000100000" => rgb <= "100001";
				when "0010000100001" => rgb <= "100001";
				when "0010000100110" => rgb <= "100001";
				when "0010000100111" => rgb <= "100001";
				when "0010000101000" => rgb <= "100001";
				when "0010000101001" => rgb <= "100001";
				when "0010000101010" => rgb <= "010000";
				when "0010000101011" => rgb <= "010000";
				when "0010000101100" => rgb <= "100001";
				when "0010000101101" => rgb <= "100001";
				when "0010000110010" => rgb <= "100001";
				when "0010000110011" => rgb <= "100001";
				when "0010000110100" => rgb <= "100001";
				when "0010000110101" => rgb <= "100001";
				when "0010000111010" => rgb <= "100001";
				when "0010000111011" => rgb <= "100001";
				when "0010000111100" => rgb <= "100001";
				when "0010000111101" => rgb <= "100001";
				when "0010001000010" => rgb <= "100001";
				when "0010001000011" => rgb <= "100001";
				when "0010001000100" => rgb <= "100001";
				when "0010001000101" => rgb <= "100001";
				when "0010001000110" => rgb <= "100001";
				when "0010001000111" => rgb <= "100001";
				when "0010001001000" => rgb <= "100100";
				when "0010001001001" => rgb <= "100100";
				when "0010010000110" => rgb <= "010000";
				when "0010010000111" => rgb <= "010000";
				when "0010010001000" => rgb <= "100001";
				when "0010010001001" => rgb <= "100001";
				when "0010010001010" => rgb <= "100001";
				when "0010010001011" => rgb <= "100001";
				when "0010010001100" => rgb <= "100001";
				when "0010010001101" => rgb <= "100001";
				when "0010010001110" => rgb <= "100001";
				when "0010010001111" => rgb <= "100001";
				when "0010010010000" => rgb <= "100001";
				when "0010010010001" => rgb <= "100001";
				when "0010010010110" => rgb <= "100001";
				when "0010010010111" => rgb <= "100001";
				when "0010010011000" => rgb <= "100001";
				when "0010010011001" => rgb <= "100001";
				when "0010010011110" => rgb <= "100001";
				when "0010010011111" => rgb <= "100001";
				when "0010010100000" => rgb <= "100001";
				when "0010010100001" => rgb <= "100001";
				when "0010010100110" => rgb <= "100001";
				when "0010010100111" => rgb <= "100100";
				when "0010010101000" => rgb <= "100100";
				when "0010010101001" => rgb <= "100100";
				when "0010010101010" => rgb <= "100100";
				when "0010010101011" => rgb <= "100001";
				when "0010010101100" => rgb <= "100001";
				when "0010010101101" => rgb <= "100001";
				when "0010010110010" => rgb <= "100001";
				when "0010010110011" => rgb <= "100100";
				when "0010010110100" => rgb <= "100100";
				when "0010010110101" => rgb <= "100001";
				when "0010010111001" => rgb <= "100001";
				when "0010010111010" => rgb <= "100100";
				when "0010010111011" => rgb <= "100001";
				when "0010010111100" => rgb <= "010000";
				when "0010010111101" => rgb <= "100001";
				when "0010011000010" => rgb <= "100100";
				when "0010011000011" => rgb <= "100001";
				when "0010011000100" => rgb <= "100001";
				when "0010011000101" => rgb <= "100001";
				when "0010011000110" => rgb <= "100100";
				when "0010011000111" => rgb <= "100100";
				when "0010011001000" => rgb <= "100100";
				when "0010011001001" => rgb <= "100001";
				when "0010100000110" => rgb <= "100100";
				when "0010100000111" => rgb <= "100100";
				when "0010100001000" => rgb <= "100100";
				when "0010100001001" => rgb <= "100001";
				when "0010100001010" => rgb <= "100001";
				when "0010100001011" => rgb <= "100001";
				when "0010100001100" => rgb <= "100001";
				when "0010100001101" => rgb <= "100100";
				when "0010100001110" => rgb <= "100100";
				when "0010100001111" => rgb <= "100100";
				when "0010100010000" => rgb <= "100100";
				when "0010100010001" => rgb <= "100001";
				when "0010100010110" => rgb <= "100001";
				when "0010100010111" => rgb <= "100001";
				when "0010100011000" => rgb <= "100001";
				when "0010100011001" => rgb <= "100001";
				when "0010100011110" => rgb <= "100001";
				when "0010100011111" => rgb <= "010000";
				when "0010100100000" => rgb <= "010000";
				when "0010100100001" => rgb <= "100001";
				when "0010100100110" => rgb <= "100001";
				when "0010100100111" => rgb <= "010000";
				when "0010100101000" => rgb <= "100001";
				when "0010100101001" => rgb <= "100001";
				when "0010100101010" => rgb <= "100001";
				when "0010100101011" => rgb <= "100001";
				when "0010100101100" => rgb <= "100001";
				when "0010100101101" => rgb <= "100001";
				when "0010100110010" => rgb <= "100001";
				when "0010100110011" => rgb <= "100001";
				when "0010100110100" => rgb <= "100100";
				when "0010100110101" => rgb <= "100001";
				when "0010100111000" => rgb <= "100001";
				when "0010100111001" => rgb <= "100001";
				when "0010100111010" => rgb <= "100001";
				when "0010100111011" => rgb <= "100001";
				when "0010100111100" => rgb <= "100001";
				when "0010101000010" => rgb <= "100001";
				when "0010101000011" => rgb <= "100001";
				when "0010101000100" => rgb <= "100001";
				when "0010101000101" => rgb <= "010000";
				when "0010101000110" => rgb <= "010000";
				when "0010101000111" => rgb <= "010000";
				when "0010101001000" => rgb <= "010000";
				when "0010101001001" => rgb <= "100001";
				when "0010110000110" => rgb <= "100001";
				when "0010110000111" => rgb <= "010000";
				when "0010110001000" => rgb <= "100100";
				when "0010110001001" => rgb <= "100100";
				when "0010110001010" => rgb <= "100001";
				when "0010110001011" => rgb <= "100001";
				when "0010110001100" => rgb <= "010000";
				when "0010110001101" => rgb <= "010000";
				when "0010110001110" => rgb <= "100001";
				when "0010110001111" => rgb <= "010000";
				when "0010110010000" => rgb <= "010000";
				when "0010110010001" => rgb <= "100001";
				when "0010110010110" => rgb <= "100001";
				when "0010110010111" => rgb <= "100100";
				when "0010110011000" => rgb <= "100001";
				when "0010110011001" => rgb <= "100001";
				when "0010110011110" => rgb <= "100001";
				when "0010110011111" => rgb <= "100100";
				when "0010110100000" => rgb <= "100001";
				when "0010110100001" => rgb <= "100001";
				when "0010110100110" => rgb <= "100001";
				when "0010110100111" => rgb <= "100001";
				when "0010110101000" => rgb <= "100001";
				when "0010110101001" => rgb <= "100001";
				when "0010110101010" => rgb <= "100001";
				when "0010110101011" => rgb <= "100001";
				when "0010110101100" => rgb <= "100001";
				when "0010110101101" => rgb <= "100001";
				when "0010110110010" => rgb <= "100001";
				when "0010110110011" => rgb <= "100001";
				when "0010110110100" => rgb <= "010000";
				when "0010110110101" => rgb <= "010000";
				when "0010110110111" => rgb <= "100001";
				when "0010110111000" => rgb <= "010000";
				when "0010110111001" => rgb <= "010000";
				when "0010110111010" => rgb <= "100001";
				when "0010110111011" => rgb <= "100001";
				when "0010111000010" => rgb <= "100001";
				when "0010111000011" => rgb <= "100001";
				when "0010111000100" => rgb <= "100001";
				when "0010111000101" => rgb <= "100001";
				when "0010111000110" => rgb <= "100001";
				when "0010111000111" => rgb <= "100001";
				when "0010111001000" => rgb <= "100001";
				when "0010111001001" => rgb <= "100001";
				when "0011000001010" => rgb <= "100001";
				when "0011000001011" => rgb <= "100001";
				when "0011000001100" => rgb <= "100001";
				when "0011000001101" => rgb <= "100001";
				when "0011000010110" => rgb <= "100001";
				when "0011000010111" => rgb <= "100001";
				when "0011000011000" => rgb <= "100001";
				when "0011000011001" => rgb <= "100001";
				when "0011000011110" => rgb <= "100001";
				when "0011000011111" => rgb <= "100001";
				when "0011000100000" => rgb <= "100001";
				when "0011000100001" => rgb <= "100001";
				when "0011000100110" => rgb <= "100100";
				when "0011000100111" => rgb <= "100100";
				when "0011000101000" => rgb <= "100100";
				when "0011000101001" => rgb <= "100001";
				when "0011000110010" => rgb <= "100001";
				when "0011000110011" => rgb <= "010000";
				when "0011000110100" => rgb <= "010000";
				when "0011000110101" => rgb <= "100001";
				when "0011000110110" => rgb <= "100001";
				when "0011000110111" => rgb <= "100100";
				when "0011000111000" => rgb <= "100100";
				when "0011000111001" => rgb <= "100100";
				when "0011000111010" => rgb <= "100001";
				when "0011001000010" => rgb <= "100001";
				when "0011001000011" => rgb <= "100001";
				when "0011001000100" => rgb <= "100100";
				when "0011001000101" => rgb <= "100001";
				when "0011010001010" => rgb <= "100001";
				when "0011010001011" => rgb <= "100001";
				when "0011010001100" => rgb <= "100001";
				when "0011010001101" => rgb <= "100001";
				when "0011010010110" => rgb <= "010000";
				when "0011010010111" => rgb <= "010000";
				when "0011010011000" => rgb <= "100001";
				when "0011010011001" => rgb <= "100001";
				when "0011010011110" => rgb <= "100001";
				when "0011010011111" => rgb <= "100100";
				when "0011010100000" => rgb <= "100001";
				when "0011010100001" => rgb <= "100001";
				when "0011010100110" => rgb <= "100001";
				when "0011010100111" => rgb <= "100001";
				when "0011010101000" => rgb <= "100001";
				when "0011010101001" => rgb <= "100001";
				when "0011010110010" => rgb <= "100001";
				when "0011010110011" => rgb <= "100001";
				when "0011010110100" => rgb <= "100001";
				when "0011010110101" => rgb <= "100001";
				when "0011010110110" => rgb <= "100001";
				when "0011010110111" => rgb <= "100001";
				when "0011010111000" => rgb <= "100001";
				when "0011010111001" => rgb <= "100001";
				when "0011011000010" => rgb <= "100001";
				when "0011011000011" => rgb <= "100001";
				when "0011011000100" => rgb <= "100001";
				when "0011011000101" => rgb <= "100001";
				when "0011100001010" => rgb <= "100001";
				when "0011100001011" => rgb <= "100001";
				when "0011100001100" => rgb <= "100001";
				when "0011100001101" => rgb <= "100001";
				when "0011100010110" => rgb <= "100001";
				when "0011100010111" => rgb <= "100001";
				when "0011100011000" => rgb <= "100001";
				when "0011100011001" => rgb <= "100001";
				when "0011100011110" => rgb <= "100001";
				when "0011100011111" => rgb <= "100001";
				when "0011100100000" => rgb <= "010000";
				when "0011100100001" => rgb <= "100001";
				when "0011100100110" => rgb <= "100001";
				when "0011100100111" => rgb <= "100100";
				when "0011100101000" => rgb <= "100001";
				when "0011100101001" => rgb <= "100001";
				when "0011100101010" => rgb <= "100001";
				when "0011100101011" => rgb <= "010000";
				when "0011100101100" => rgb <= "010000";
				when "0011100101101" => rgb <= "010000";
				when "0011100110010" => rgb <= "100001";
				when "0011100110011" => rgb <= "100001";
				when "0011100110100" => rgb <= "100001";
				when "0011100110101" => rgb <= "100001";
				when "0011100110110" => rgb <= "100001";
				when "0011100110111" => rgb <= "100001";
				when "0011100111000" => rgb <= "100001";
				when "0011101000010" => rgb <= "100001";
				when "0011101000011" => rgb <= "100001";
				when "0011101000100" => rgb <= "100001";
				when "0011101000101" => rgb <= "100001";
				when "0011101000110" => rgb <= "100001";
				when "0011101000111" => rgb <= "100001";
				when "0011101001000" => rgb <= "100001";
				when "0011101001001" => rgb <= "100001";
				when "0011110001010" => rgb <= "100001";
				when "0011110001011" => rgb <= "100001";
				when "0011110001100" => rgb <= "100001";
				when "0011110001101" => rgb <= "100001";
				when "0011110010110" => rgb <= "100001";
				when "0011110010111" => rgb <= "100100";
				when "0011110011000" => rgb <= "100100";
				when "0011110011001" => rgb <= "100001";
				when "0011110011110" => rgb <= "010000";
				when "0011110011111" => rgb <= "010000";
				when "0011110100000" => rgb <= "100001";
				when "0011110100001" => rgb <= "100100";
				when "0011110100110" => rgb <= "100001";
				when "0011110100111" => rgb <= "100001";
				when "0011110101000" => rgb <= "100001";
				when "0011110101001" => rgb <= "100001";
				when "0011110101010" => rgb <= "100100";
				when "0011110101011" => rgb <= "100100";
				when "0011110101100" => rgb <= "100100";
				when "0011110101101" => rgb <= "100001";
				when "0011110110010" => rgb <= "100001";
				when "0011110110011" => rgb <= "100001";
				when "0011110110100" => rgb <= "100001";
				when "0011110110101" => rgb <= "010000";
				when "0011110110110" => rgb <= "010000";
				when "0011110110111" => rgb <= "010000";
				when "0011110111000" => rgb <= "100001";
				when "0011111000010" => rgb <= "100001";
				when "0011111000011" => rgb <= "100001";
				when "0011111000100" => rgb <= "100001";
				when "0011111000101" => rgb <= "100001";
				when "0011111000110" => rgb <= "010000";
				when "0011111000111" => rgb <= "100001";
				when "0011111001000" => rgb <= "100100";
				when "0011111001001" => rgb <= "100100";
				when "0100000001010" => rgb <= "010000";
				when "0100000001011" => rgb <= "100001";
				when "0100000001100" => rgb <= "100001";
				when "0100000001101" => rgb <= "100001";
				when "0100000010110" => rgb <= "100001";
				when "0100000010111" => rgb <= "100001";
				when "0100000011000" => rgb <= "100100";
				when "0100000011001" => rgb <= "100001";
				when "0100000011110" => rgb <= "100001";
				when "0100000011111" => rgb <= "100001";
				when "0100000100000" => rgb <= "100001";
				when "0100000100001" => rgb <= "100001";
				when "0100000101010" => rgb <= "100001";
				when "0100000101011" => rgb <= "100001";
				when "0100000101100" => rgb <= "100100";
				when "0100000101101" => rgb <= "100100";
				when "0100000110010" => rgb <= "100001";
				when "0100000110011" => rgb <= "100100";
				when "0100000110100" => rgb <= "100100";
				when "0100000110101" => rgb <= "100100";
				when "0100000110110" => rgb <= "100100";
				when "0100000110111" => rgb <= "100100";
				when "0100000111000" => rgb <= "100001";
				when "0100000111001" => rgb <= "100001";
				when "0100001000110" => rgb <= "100001";
				when "0100001000111" => rgb <= "100001";
				when "0100001001000" => rgb <= "010000";
				when "0100001001001" => rgb <= "100001";
				when "0100010001010" => rgb <= "100001";
				when "0100010001011" => rgb <= "100001";
				when "0100010001100" => rgb <= "100001";
				when "0100010001101" => rgb <= "100001";
				when "0100010010110" => rgb <= "100001";
				when "0100010010111" => rgb <= "100001";
				when "0100010011000" => rgb <= "100001";
				when "0100010011001" => rgb <= "100001";
				when "0100010011110" => rgb <= "100001";
				when "0100010011111" => rgb <= "100001";
				when "0100010100000" => rgb <= "100001";
				when "0100010100001" => rgb <= "100001";
				when "0100010101010" => rgb <= "010000";
				when "0100010101011" => rgb <= "010000";
				when "0100010101100" => rgb <= "100001";
				when "0100010101101" => rgb <= "100001";
				when "0100010110010" => rgb <= "100001";
				when "0100010110011" => rgb <= "100001";
				when "0100010110100" => rgb <= "100001";
				when "0100010110101" => rgb <= "100001";
				when "0100010110110" => rgb <= "100001";
				when "0100010110111" => rgb <= "100100";
				when "0100010111000" => rgb <= "100100";
				when "0100010111001" => rgb <= "100100";
				when "0100010111010" => rgb <= "010000";
				when "0100011000110" => rgb <= "100001";
				when "0100011000111" => rgb <= "100100";
				when "0100011001000" => rgb <= "100001";
				when "0100011001001" => rgb <= "100001";
				when "0100100001010" => rgb <= "100001";
				when "0100100001011" => rgb <= "100001";
				when "0100100001100" => rgb <= "100001";
				when "0100100001101" => rgb <= "100001";
				when "0100100010110" => rgb <= "100001";
				when "0100100010111" => rgb <= "010000";
				when "0100100011000" => rgb <= "010000";
				when "0100100011001" => rgb <= "100001";
				when "0100100011010" => rgb <= "100001";
				when "0100100011011" => rgb <= "100100";
				when "0100100011100" => rgb <= "100100";
				when "0100100011101" => rgb <= "100100";
				when "0100100011110" => rgb <= "100001";
				when "0100100011111" => rgb <= "010000";
				when "0100100100000" => rgb <= "010000";
				when "0100100100001" => rgb <= "100001";
				when "0100100100110" => rgb <= "100001";
				when "0100100100111" => rgb <= "100100";
				when "0100100101000" => rgb <= "100001";
				when "0100100101001" => rgb <= "100001";
				when "0100100101010" => rgb <= "100001";
				when "0100100101011" => rgb <= "100001";
				when "0100100101100" => rgb <= "100001";
				when "0100100101101" => rgb <= "100001";
				when "0100100110010" => rgb <= "100001";
				when "0100100110011" => rgb <= "100001";
				when "0100100110100" => rgb <= "100001";
				when "0100100110101" => rgb <= "100001";
				when "0100100110111" => rgb <= "100001";
				when "0100100111000" => rgb <= "100001";
				when "0100100111001" => rgb <= "010000";
				when "0100100111010" => rgb <= "010000";
				when "0100100111011" => rgb <= "100001";
				when "0100101000010" => rgb <= "100001";
				when "0100101000011" => rgb <= "100001";
				when "0100101000100" => rgb <= "100001";
				when "0100101000101" => rgb <= "100001";
				when "0100101000110" => rgb <= "010000";
				when "0100101000111" => rgb <= "100001";
				when "0100101001000" => rgb <= "100001";
				when "0100101001001" => rgb <= "100001";
				when "0100110001010" => rgb <= "100001";
				when "0100110001011" => rgb <= "100001";
				when "0100110001100" => rgb <= "010000";
				when "0100110001101" => rgb <= "100001";
				when "0100110010110" => rgb <= "100001";
				when "0100110010111" => rgb <= "100001";
				when "0100110011000" => rgb <= "100100";
				when "0100110011001" => rgb <= "100001";
				when "0100110011010" => rgb <= "010000";
				when "0100110011011" => rgb <= "010000";
				when "0100110011100" => rgb <= "010000";
				when "0100110011101" => rgb <= "100001";
				when "0100110011110" => rgb <= "100001";
				when "0100110011111" => rgb <= "100001";
				when "0100110100000" => rgb <= "100001";
				when "0100110100001" => rgb <= "100001";
				when "0100110100110" => rgb <= "010000";
				when "0100110100111" => rgb <= "100001";
				when "0100110101000" => rgb <= "100001";
				when "0100110101001" => rgb <= "100001";
				when "0100110101010" => rgb <= "100001";
				when "0100110101011" => rgb <= "100001";
				when "0100110101100" => rgb <= "100001";
				when "0100110101101" => rgb <= "100001";
				when "0100110110010" => rgb <= "100001";
				when "0100110110011" => rgb <= "100100";
				when "0100110110100" => rgb <= "100001";
				when "0100110110101" => rgb <= "100001";
				when "0100110111000" => rgb <= "100001";
				when "0100110111001" => rgb <= "100001";
				when "0100110111010" => rgb <= "100001";
				when "0100110111011" => rgb <= "100001";
				when "0100110111100" => rgb <= "100001";
				when "0100111000010" => rgb <= "100001";
				when "0100111000011" => rgb <= "100001";
				when "0100111000100" => rgb <= "100001";
				when "0100111000101" => rgb <= "100001";
				when "0100111000110" => rgb <= "100001";
				when "0100111000111" => rgb <= "100100";
				when "0100111001000" => rgb <= "100100";
				when "0100111001001" => rgb <= "100100";
				when "0101000001010" => rgb <= "100001";
				when "0101000001011" => rgb <= "100100";
				when "0101000001100" => rgb <= "100001";
				when "0101000001101" => rgb <= "010000";
				when "0101000011000" => rgb <= "100001";
				when "0101000011001" => rgb <= "100001";
				when "0101000011010" => rgb <= "100001";
				when "0101000011011" => rgb <= "100001";
				when "0101000011100" => rgb <= "100001";
				when "0101000011101" => rgb <= "100100";
				when "0101000011110" => rgb <= "100100";
				when "0101000011111" => rgb <= "100001";
				when "0101000100110" => rgb <= "100001";
				when "0101000100111" => rgb <= "001011";
				when "0101000101000" => rgb <= "100001";
				when "0101000101001" => rgb <= "010000";
				when "0101000101010" => rgb <= "100001";
				when "0101000101011" => rgb <= "100100";
				when "0101000101100" => rgb <= "100100";
				when "0101000101101" => rgb <= "100001";
				when "0101000110010" => rgb <= "100001";
				when "0101000110011" => rgb <= "100001";
				when "0101000110100" => rgb <= "100100";
				when "0101000110101" => rgb <= "100001";
				when "0101000111001" => rgb <= "100001";
				when "0101000111010" => rgb <= "100001";
				when "0101000111011" => rgb <= "100100";
				when "0101000111100" => rgb <= "100100";
				when "0101000111101" => rgb <= "100001";
				when "0101001000010" => rgb <= "100001";
				when "0101001000011" => rgb <= "100001";
				when "0101001000100" => rgb <= "100001";
				when "0101001000101" => rgb <= "100100";
				when "0101001000110" => rgb <= "100001";
				when "0101001000111" => rgb <= "100001";
				when "0101001001000" => rgb <= "100100";
				when "0101001001001" => rgb <= "100001";
				when "0101010001010" => rgb <= "010000";
				when "0101010001011" => rgb <= "100001";
				when "0101010001100" => rgb <= "100001";
				when "0101010001101" => rgb <= "100001";
				when "0101010011000" => rgb <= "100100";
				when "0101010011001" => rgb <= "100001";
				when "0101010011010" => rgb <= "100001";
				when "0101010011011" => rgb <= "100001";
				when "0101010011100" => rgb <= "010000";
				when "0101010011101" => rgb <= "100001";
				when "0101010011110" => rgb <= "100001";
				when "0101010011111" => rgb <= "100001";
				when "0101010100110" => rgb <= "100001";
				when "0101010100111" => rgb <= "001011";
				when "0101010101000" => rgb <= "100001";
				when "0101010101001" => rgb <= "100001";
				when "0101010101010" => rgb <= "010000";
				when "0101010101011" => rgb <= "010000";
				when "0101010101100" => rgb <= "010000";
				when "0101010101101" => rgb <= "100001";
				when "0101010110010" => rgb <= "100001";
				when "0101010110011" => rgb <= "100001";
				when "0101010110100" => rgb <= "100001";
				when "0101010110101" => rgb <= "100001";
				when "0101010111010" => rgb <= "010000";
				when "0101010111011" => rgb <= "010000";
				when "0101010111100" => rgb <= "100001";
				when "0101010111101" => rgb <= "100001";
				when "0101011000010" => rgb <= "010000";
				when "0101011000011" => rgb <= "100001";
				when "0101011000100" => rgb <= "100001";
				when "0101011000101" => rgb <= "100001";
				when "0101011000110" => rgb <= "100001";
				when "0101011000111" => rgb <= "100001";
				when "0101011001000" => rgb <= "100001";
				when "0101011001001" => rgb <= "100001";
				when "0110100100100" => rgb <= "111111";
				when "0110100100101" => rgb <= "111111";
				when "0110100100110" => rgb <= "111111";
				when "0110100100111" => rgb <= "111111";
				when "0110100101000" => rgb <= "111111";
				when "0110100101001" => rgb <= "111111";
				when "0110100101010" => rgb <= "111111";
				when "0110100101011" => rgb <= "111111";
				when "0110100101100" => rgb <= "111111";
				when "0110100101101" => rgb <= "111111";
				when "0110110100100" => rgb <= "111111";
				when "0110110100101" => rgb <= "111111";
				when "0110110100110" => rgb <= "111111";
				when "0110110100111" => rgb <= "111111";
				when "0110110101000" => rgb <= "111111";
				when "0110110101001" => rgb <= "111111";
				when "0110110101010" => rgb <= "111111";
				when "0110110101011" => rgb <= "111111";
				when "0110110101100" => rgb <= "111111";
				when "0110110101101" => rgb <= "111111";
				when "0111000011110" => rgb <= "111111";
				when "0111000011111" => rgb <= "111111";
				when "0111000100000" => rgb <= "111111";
				when "0111000100001" => rgb <= "111111";
				when "0111000100010" => rgb <= "111111";
				when "0111000100011" => rgb <= "111111";
				when "0111000100100" => rgb <= "111111";
				when "0111000100101" => rgb <= "111111";
				when "0111000100110" => rgb <= "111111";
				when "0111000100111" => rgb <= "111111";
				when "0111000101000" => rgb <= "111111";
				when "0111000101001" => rgb <= "111111";
				when "0111000101010" => rgb <= "111111";
				when "0111000101011" => rgb <= "111111";
				when "0111000101100" => rgb <= "111111";
				when "0111000101101" => rgb <= "111111";
				when "0111000101110" => rgb <= "111111";
				when "0111000101111" => rgb <= "111111";
				when "0111010011110" => rgb <= "111111";
				when "0111010011111" => rgb <= "111111";
				when "0111010100000" => rgb <= "111111";
				when "0111010100001" => rgb <= "111111";
				when "0111010100010" => rgb <= "111111";
				when "0111010100011" => rgb <= "111111";
				when "0111010100100" => rgb <= "111111";
				when "0111010100101" => rgb <= "111111";
				when "0111010100110" => rgb <= "111111";
				when "0111010100111" => rgb <= "111111";
				when "0111010101000" => rgb <= "111111";
				when "0111010101001" => rgb <= "111111";
				when "0111010101010" => rgb <= "111111";
				when "0111010101011" => rgb <= "111111";
				when "0111010101100" => rgb <= "111111";
				when "0111010101101" => rgb <= "111111";
				when "0111010101110" => rgb <= "111111";
				when "0111010101111" => rgb <= "111111";
				when "0111100011100" => rgb <= "111111";
				when "0111100011101" => rgb <= "111111";
				when "0111100011110" => rgb <= "111111";
				when "0111100011111" => rgb <= "111111";
				when "0111100100000" => rgb <= "111111";
				when "0111100100001" => rgb <= "111111";
				when "0111100100010" => rgb <= "111111";
				when "0111100100011" => rgb <= "111111";
				when "0111100100100" => rgb <= "111111";
				when "0111100100101" => rgb <= "111111";
				when "0111100100110" => rgb <= "111111";
				when "0111100100111" => rgb <= "111111";
				when "0111100101000" => rgb <= "111111";
				when "0111100101001" => rgb <= "111111";
				when "0111100101010" => rgb <= "111111";
				when "0111100101011" => rgb <= "111111";
				when "0111100101100" => rgb <= "111111";
				when "0111100101101" => rgb <= "111111";
				when "0111100101110" => rgb <= "111111";
				when "0111100101111" => rgb <= "111111";
				when "0111110011100" => rgb <= "111111";
				when "0111110011101" => rgb <= "111111";
				when "0111110011110" => rgb <= "111111";
				when "0111110011111" => rgb <= "111111";
				when "0111110100000" => rgb <= "111111";
				when "0111110100001" => rgb <= "111111";
				when "0111110100010" => rgb <= "111111";
				when "0111110100011" => rgb <= "111111";
				when "0111110100100" => rgb <= "111111";
				when "0111110100101" => rgb <= "111111";
				when "0111110100110" => rgb <= "111111";
				when "0111110100111" => rgb <= "111111";
				when "0111110101000" => rgb <= "111111";
				when "0111110101001" => rgb <= "111111";
				when "0111110101010" => rgb <= "111111";
				when "0111110101011" => rgb <= "111111";
				when "0111110101100" => rgb <= "111111";
				when "0111110101101" => rgb <= "111111";
				when "0111110101110" => rgb <= "111111";
				when "0111110101111" => rgb <= "111111";
				when "1000000011010" => rgb <= "111111";
				when "1000000011011" => rgb <= "111111";
				when "1000000011100" => rgb <= "111111";
				when "1000000011101" => rgb <= "111111";
				when "1000000011110" => rgb <= "111111";
				when "1000000011111" => rgb <= "111111";
				when "1000000100000" => rgb <= "111111";
				when "1000000100001" => rgb <= "111111";
				when "1000000100010" => rgb <= "111111";
				when "1000000100011" => rgb <= "111111";
				when "1000000100100" => rgb <= "111111";
				when "1000000100101" => rgb <= "111111";
				when "1000000100110" => rgb <= "111111";
				when "1000000100111" => rgb <= "111111";
				when "1000000101000" => rgb <= "111111";
				when "1000000101001" => rgb <= "111111";
				when "1000000101100" => rgb <= "111111";
				when "1000000101101" => rgb <= "111111";
				when "1000000101110" => rgb <= "111111";
				when "1000000101111" => rgb <= "111111";
				when "1000010011010" => rgb <= "111111";
				when "1000010011011" => rgb <= "111111";
				when "1000010011100" => rgb <= "111111";
				when "1000010011101" => rgb <= "111111";
				when "1000010011110" => rgb <= "111111";
				when "1000010011111" => rgb <= "111111";
				when "1000010100000" => rgb <= "111111";
				when "1000010100001" => rgb <= "111111";
				when "1000010100010" => rgb <= "111111";
				when "1000010100011" => rgb <= "111111";
				when "1000010100100" => rgb <= "111111";
				when "1000010100101" => rgb <= "111111";
				when "1000010100110" => rgb <= "111111";
				when "1000010100111" => rgb <= "111111";
				when "1000010101000" => rgb <= "111111";
				when "1000010101001" => rgb <= "111111";
				when "1000010101100" => rgb <= "111111";
				when "1000010101101" => rgb <= "111111";
				when "1000010101110" => rgb <= "111111";
				when "1000010101111" => rgb <= "111111";
				when "1000100011000" => rgb <= "111111";
				when "1000100011001" => rgb <= "111111";
				when "1000100011010" => rgb <= "111111";
				when "1000100011011" => rgb <= "111111";
				when "1000100011100" => rgb <= "111111";
				when "1000100011101" => rgb <= "111111";
				when "1000100011110" => rgb <= "111111";
				when "1000100011111" => rgb <= "111111";
				when "1000100100000" => rgb <= "111111";
				when "1000100100001" => rgb <= "111111";
				when "1000100100010" => rgb <= "111111";
				when "1000100100011" => rgb <= "111111";
				when "1000100100100" => rgb <= "111111";
				when "1000100100101" => rgb <= "111111";
				when "1000100100110" => rgb <= "111111";
				when "1000100100111" => rgb <= "111111";
				when "1000100101000" => rgb <= "111111";
				when "1000100101001" => rgb <= "111111";
				when "1000100101010" => rgb <= "111111";
				when "1000100101011" => rgb <= "111111";
				when "1000100101100" => rgb <= "111111";
				when "1000100101101" => rgb <= "111111";
				when "1000100101110" => rgb <= "111111";
				when "1000100101111" => rgb <= "111111";
				when "1000110011000" => rgb <= "111111";
				when "1000110011001" => rgb <= "111111";
				when "1000110011010" => rgb <= "111111";
				when "1000110011011" => rgb <= "111111";
				when "1000110011100" => rgb <= "111111";
				when "1000110011101" => rgb <= "111111";
				when "1000110011110" => rgb <= "111111";
				when "1000110011111" => rgb <= "111111";
				when "1000110100000" => rgb <= "111111";
				when "1000110100001" => rgb <= "111111";
				when "1000110100010" => rgb <= "111111";
				when "1000110100011" => rgb <= "111111";
				when "1000110100100" => rgb <= "111111";
				when "1000110100101" => rgb <= "111111";
				when "1000110100110" => rgb <= "111111";
				when "1000110100111" => rgb <= "111111";
				when "1000110101000" => rgb <= "111111";
				when "1000110101001" => rgb <= "111111";
				when "1000110101010" => rgb <= "111111";
				when "1000110101011" => rgb <= "111111";
				when "1000110101100" => rgb <= "111111";
				when "1000110101101" => rgb <= "111111";
				when "1000110101110" => rgb <= "111111";
				when "1000110101111" => rgb <= "111111";
				when "1001000011010" => rgb <= "111111";
				when "1001000011011" => rgb <= "111111";
				when "1001000011100" => rgb <= "111111";
				when "1001000011101" => rgb <= "111111";
				when "1001000011110" => rgb <= "111111";
				when "1001000011111" => rgb <= "111111";
				when "1001000100000" => rgb <= "111111";
				when "1001000100001" => rgb <= "111111";
				when "1001000100010" => rgb <= "111111";
				when "1001000100011" => rgb <= "111111";
				when "1001000100100" => rgb <= "111111";
				when "1001000100101" => rgb <= "111111";
				when "1001000100110" => rgb <= "111111";
				when "1001000100111" => rgb <= "111111";
				when "1001000101000" => rgb <= "111111";
				when "1001000101001" => rgb <= "111111";
				when "1001000101010" => rgb <= "111111";
				when "1001000101011" => rgb <= "111111";
				when "1001000101100" => rgb <= "111111";
				when "1001000101101" => rgb <= "111111";
				when "1001000101110" => rgb <= "111111";
				when "1001000101111" => rgb <= "111111";
				when "1001010011010" => rgb <= "111111";
				when "1001010011011" => rgb <= "111111";
				when "1001010011100" => rgb <= "111111";
				when "1001010011101" => rgb <= "111111";
				when "1001010011110" => rgb <= "111111";
				when "1001010011111" => rgb <= "111111";
				when "1001010100000" => rgb <= "111111";
				when "1001010100001" => rgb <= "111111";
				when "1001010100010" => rgb <= "111111";
				when "1001010100011" => rgb <= "111111";
				when "1001010100100" => rgb <= "111111";
				when "1001010100101" => rgb <= "111111";
				when "1001010100110" => rgb <= "111111";
				when "1001010100111" => rgb <= "111111";
				when "1001010101000" => rgb <= "111111";
				when "1001010101001" => rgb <= "111111";
				when "1001010101010" => rgb <= "111111";
				when "1001010101011" => rgb <= "111111";
				when "1001010101100" => rgb <= "111111";
				when "1001010101101" => rgb <= "111111";
				when "1001010101110" => rgb <= "111111";
				when "1001010101111" => rgb <= "111111";
				when "1001100011010" => rgb <= "111111";
				when "1001100011011" => rgb <= "111111";
				when "1001100011100" => rgb <= "111111";
				when "1001100011101" => rgb <= "111111";
				when "1001100011110" => rgb <= "111111";
				when "1001100011111" => rgb <= "111111";
				when "1001100100000" => rgb <= "111111";
				when "1001100100001" => rgb <= "111111";
				when "1001100100010" => rgb <= "111111";
				when "1001100100011" => rgb <= "111111";
				when "1001100100100" => rgb <= "111111";
				when "1001100100101" => rgb <= "111111";
				when "1001100100110" => rgb <= "111111";
				when "1001100100111" => rgb <= "111111";
				when "1001100101000" => rgb <= "111111";
				when "1001100101001" => rgb <= "111111";
				when "1001100101010" => rgb <= "111111";
				when "1001100101011" => rgb <= "111111";
				when "1001100101100" => rgb <= "111111";
				when "1001100101101" => rgb <= "111111";
				when "1001100101110" => rgb <= "111111";
				when "1001100101111" => rgb <= "111111";
				when "1001110011010" => rgb <= "111111";
				when "1001110011011" => rgb <= "111111";
				when "1001110011100" => rgb <= "111111";
				when "1001110011101" => rgb <= "111111";
				when "1001110011110" => rgb <= "111111";
				when "1001110011111" => rgb <= "111111";
				when "1001110100000" => rgb <= "111111";
				when "1001110100001" => rgb <= "111111";
				when "1001110100010" => rgb <= "111111";
				when "1001110100011" => rgb <= "111111";
				when "1001110100100" => rgb <= "111111";
				when "1001110100101" => rgb <= "111111";
				when "1001110100110" => rgb <= "111111";
				when "1001110100111" => rgb <= "111111";
				when "1001110101000" => rgb <= "111111";
				when "1001110101001" => rgb <= "111111";
				when "1001110101010" => rgb <= "111111";
				when "1001110101011" => rgb <= "111111";
				when "1001110101100" => rgb <= "111111";
				when "1001110101101" => rgb <= "111111";
				when "1001110101110" => rgb <= "111111";
				when "1001110101111" => rgb <= "111111";
				when "1010000011010" => rgb <= "111111";
				when "1010000011011" => rgb <= "111111";
				when "1010000011100" => rgb <= "111111";
				when "1010000011101" => rgb <= "111111";
				when "1010000011110" => rgb <= "111111";
				when "1010000011111" => rgb <= "111111";
				when "1010000100100" => rgb <= "111111";
				when "1010000100101" => rgb <= "111111";
				when "1010000100110" => rgb <= "111111";
				when "1010000100111" => rgb <= "111111";
				when "1010000101000" => rgb <= "111111";
				when "1010000101001" => rgb <= "111111";
				when "1010000101100" => rgb <= "111111";
				when "1010000101101" => rgb <= "111111";
				when "1010000101110" => rgb <= "111111";
				when "1010000101111" => rgb <= "111111";
				when "1010000110000" => rgb <= "111111";
				when "1010000110001" => rgb <= "111111";
				when "1010010011010" => rgb <= "111111";
				when "1010010011011" => rgb <= "111111";
				when "1010010011100" => rgb <= "111111";
				when "1010010011101" => rgb <= "111111";
				when "1010010011110" => rgb <= "111111";
				when "1010010011111" => rgb <= "111111";
				when "1010010100100" => rgb <= "111111";
				when "1010010100101" => rgb <= "111111";
				when "1010010100110" => rgb <= "111111";
				when "1010010100111" => rgb <= "111111";
				when "1010010101000" => rgb <= "111111";
				when "1010010101001" => rgb <= "111111";
				when "1010010101100" => rgb <= "111111";
				when "1010010101101" => rgb <= "111111";
				when "1010010101110" => rgb <= "111111";
				when "1010010101111" => rgb <= "111111";
				when "1010010110000" => rgb <= "111111";
				when "1010010110001" => rgb <= "111111";
				when "1010100011010" => rgb <= "111111";
				when "1010100011011" => rgb <= "111111";
				when "1010100011100" => rgb <= "111111";
				when "1010100011101" => rgb <= "111111";
				when "1010100011110" => rgb <= "111111";
				when "1010100011111" => rgb <= "111111";
				when "1010100100100" => rgb <= "111111";
				when "1010100100101" => rgb <= "111111";
				when "1010100100110" => rgb <= "111111";
				when "1010100100111" => rgb <= "111111";
				when "1010100101000" => rgb <= "111111";
				when "1010100101001" => rgb <= "111111";
				when "1010100110000" => rgb <= "111111";
				when "1010100110001" => rgb <= "111111";
				when "1010100110010" => rgb <= "111111";
				when "1010100110011" => rgb <= "111111";
				when "1010110011010" => rgb <= "111111";
				when "1010110011011" => rgb <= "111111";
				when "1010110011100" => rgb <= "111111";
				when "1010110011101" => rgb <= "111111";
				when "1010110011110" => rgb <= "111111";
				when "1010110011111" => rgb <= "111111";
				when "1010110100100" => rgb <= "111111";
				when "1010110100101" => rgb <= "111111";
				when "1010110100110" => rgb <= "111111";
				when "1010110100111" => rgb <= "111111";
				when "1010110101000" => rgb <= "111111";
				when "1010110101001" => rgb <= "111111";
				when "1010110110000" => rgb <= "111111";
				when "1010110110001" => rgb <= "111111";
				when "1010110110010" => rgb <= "111111";
				when "1010110110011" => rgb <= "111111";
				when "1011000011010" => rgb <= "111111";
				when "1011000011011" => rgb <= "111111";
				when "1011000011100" => rgb <= "111111";
				when "1011000011101" => rgb <= "111111";
				when "1011000011110" => rgb <= "111111";
				when "1011000011111" => rgb <= "111111";
				when "1011000100100" => rgb <= "111111";
				when "1011000100101" => rgb <= "111111";
				when "1011000100110" => rgb <= "111111";
				when "1011000100111" => rgb <= "111111";
				when "1011000101000" => rgb <= "111111";
				when "1011000101001" => rgb <= "111111";
				when "1011010011010" => rgb <= "111111";
				when "1011010011011" => rgb <= "111111";
				when "1011010011100" => rgb <= "111111";
				when "1011010011101" => rgb <= "111111";
				when "1011010011110" => rgb <= "111111";
				when "1011010011111" => rgb <= "111111";
				when "1011010100100" => rgb <= "111111";
				when "1011010100101" => rgb <= "111111";
				when "1011010100110" => rgb <= "111111";
				when "1011010100111" => rgb <= "111111";
				when "1011010101000" => rgb <= "111111";
				when "1011010101001" => rgb <= "111111";
				when "1100000011101" => rgb <= "111111";
				when "1100000011110" => rgb <= "111111";
				when "1100000011111" => rgb <= "111111";
				when "1100000100000" => rgb <= "111111";
				when "1100000100001" => rgb <= "111111";
				when "1100000100010" => rgb <= "111111";
				when "1100000100011" => rgb <= "111111";
				when "1100000100100" => rgb <= "111111";
				when "1100000100101" => rgb <= "111111";
				when "1100000100110" => rgb <= "111111";
				when "1100000100111" => rgb <= "111111";
				when "1100000101000" => rgb <= "111111";
				when "1100000101001" => rgb <= "111111";
				when "1100000101010" => rgb <= "111111";
				when "1100000101011" => rgb <= "111111";
				when "1100000101100" => rgb <= "111111";
				when "1100000101101" => rgb <= "111111";
				when "1100000101110" => rgb <= "111111";
				when "1100010011100" => rgb <= "001011";
				when "1100010011101" => rgb <= "001011";
				when "1100010011110" => rgb <= "001011";
				when "1100010011111" => rgb <= "001011";
				when "1100010100000" => rgb <= "001011";
				when "1100010100001" => rgb <= "001011";
				when "1100010100010" => rgb <= "001011";
				when "1100010100011" => rgb <= "001011";
				when "1100010100100" => rgb <= "001011";
				when "1100010100101" => rgb <= "001011";
				when "1100010100110" => rgb <= "001011";
				when "1100010100111" => rgb <= "001011";
				when "1100010101000" => rgb <= "001011";
				when "1100010101001" => rgb <= "001011";
				when "1100010101010" => rgb <= "001011";
				when "1100010101011" => rgb <= "001011";
				when "1100010101100" => rgb <= "001011";
				when "1100010101101" => rgb <= "001011";
				when "1100010101110" => rgb <= "001011";
				when "1100010101111" => rgb <= "001011";
				when "1100100011011" => rgb <= "111111";
				when "1100100011100" => rgb <= "001011";
				when "1100100011101" => rgb <= "001011";
				when "1100100011110" => rgb <= "001011";
				when "1100100011111" => rgb <= "111111";
				when "1100100100000" => rgb <= "111111";
				when "1100100100001" => rgb <= "111111";
				when "1100100100010" => rgb <= "001011";
				when "1100100100011" => rgb <= "111111";
				when "1100100100100" => rgb <= "001011";
				when "1100100100101" => rgb <= "001011";
				when "1100100100110" => rgb <= "111111";
				when "1100100100111" => rgb <= "111111";
				when "1100100101000" => rgb <= "111111";
				when "1100100101001" => rgb <= "001011";
				when "1100100101010" => rgb <= "111111";
				when "1100100101011" => rgb <= "001011";
				when "1100100101100" => rgb <= "111111";
				when "1100100101101" => rgb <= "001011";
				when "1100100101110" => rgb <= "001011";
				when "1100100101111" => rgb <= "001011";
				when "1100100110000" => rgb <= "111111";
				when "1100110011011" => rgb <= "111111";
				when "1100110011100" => rgb <= "001011";
				when "1100110011101" => rgb <= "001011";
				when "1100110011110" => rgb <= "001011";
				when "1100110011111" => rgb <= "111111";
				when "1100110100000" => rgb <= "001011";
				when "1100110100001" => rgb <= "111111";
				when "1100110100010" => rgb <= "001011";
				when "1100110100011" => rgb <= "111111";
				when "1100110100100" => rgb <= "001011";
				when "1100110100101" => rgb <= "001011";
				when "1100110100110" => rgb <= "111111";
				when "1100110100111" => rgb <= "001011";
				when "1100110101000" => rgb <= "111111";
				when "1100110101001" => rgb <= "001011";
				when "1100110101010" => rgb <= "111111";
				when "1100110101011" => rgb <= "001011";
				when "1100110101100" => rgb <= "111111";
				when "1100110101101" => rgb <= "001011";
				when "1100110101110" => rgb <= "001011";
				when "1100110101111" => rgb <= "001011";
				when "1100110110000" => rgb <= "111111";
				when "1101000011011" => rgb <= "111111";
				when "1101000011100" => rgb <= "001011";
				when "1101000011101" => rgb <= "001011";
				when "1101000011110" => rgb <= "001011";
				when "1101000011111" => rgb <= "111111";
				when "1101000100000" => rgb <= "111111";
				when "1101000100001" => rgb <= "111111";
				when "1101000100010" => rgb <= "001011";
				when "1101000100011" => rgb <= "111111";
				when "1101000100100" => rgb <= "001011";
				when "1101000100101" => rgb <= "001011";
				when "1101000100110" => rgb <= "111111";
				when "1101000100111" => rgb <= "111111";
				when "1101000101000" => rgb <= "111111";
				when "1101000101001" => rgb <= "001011";
				when "1101000101010" => rgb <= "001011";
				when "1101000101011" => rgb <= "111111";
				when "1101000101100" => rgb <= "001011";
				when "1101000101101" => rgb <= "001011";
				when "1101000101110" => rgb <= "001011";
				when "1101000101111" => rgb <= "001011";
				when "1101000110000" => rgb <= "111111";
				when "1101010011011" => rgb <= "111111";
				when "1101010011100" => rgb <= "001011";
				when "1101010011101" => rgb <= "001011";
				when "1101010011110" => rgb <= "001011";
				when "1101010011111" => rgb <= "111111";
				when "1101010100000" => rgb <= "001011";
				when "1101010100001" => rgb <= "001011";
				when "1101010100010" => rgb <= "001011";
				when "1101010100011" => rgb <= "111111";
				when "1101010100100" => rgb <= "111111";
				when "1101010100101" => rgb <= "001011";
				when "1101010100110" => rgb <= "111111";
				when "1101010100111" => rgb <= "001011";
				when "1101010101000" => rgb <= "111111";
				when "1101010101001" => rgb <= "001011";
				when "1101010101010" => rgb <= "001011";
				when "1101010101011" => rgb <= "111111";
				when "1101010101100" => rgb <= "001011";
				when "1101010101101" => rgb <= "001011";
				when "1101010101110" => rgb <= "001011";
				when "1101010101111" => rgb <= "001011";
				when "1101010110000" => rgb <= "111111";
				when "1101100011100" => rgb <= "000110";
				when "1101100011101" => rgb <= "001011";
				when "1101100011110" => rgb <= "001011";
				when "1101100011111" => rgb <= "001011";
				when "1101100100000" => rgb <= "001011";
				when "1101100100001" => rgb <= "001011";
				when "1101100100010" => rgb <= "001011";
				when "1101100100011" => rgb <= "001011";
				when "1101100100100" => rgb <= "001011";
				when "1101100100101" => rgb <= "001011";
				when "1101100100110" => rgb <= "001011";
				when "1101100100111" => rgb <= "001011";
				when "1101100101000" => rgb <= "001011";
				when "1101100101001" => rgb <= "001011";
				when "1101100101010" => rgb <= "001011";
				when "1101100101011" => rgb <= "001011";
				when "1101100101100" => rgb <= "001011";
				when "1101100101101" => rgb <= "001011";
				when "1101100101110" => rgb <= "001011";
				when "1101100101111" => rgb <= "000110";
				when "1101110011100" => rgb <= "111111";
				when "1101110011101" => rgb <= "000110";
				when "1101110011110" => rgb <= "000110";
				when "1101110011111" => rgb <= "000110";
				when "1101110100000" => rgb <= "000110";
				when "1101110100001" => rgb <= "000110";
				when "1101110100010" => rgb <= "000110";
				when "1101110100011" => rgb <= "000110";
				when "1101110100100" => rgb <= "000110";
				when "1101110100101" => rgb <= "000110";
				when "1101110100110" => rgb <= "000110";
				when "1101110100111" => rgb <= "000110";
				when "1101110101000" => rgb <= "000110";
				when "1101110101001" => rgb <= "000110";
				when "1101110101010" => rgb <= "000110";
				when "1101110101011" => rgb <= "000110";
				when "1101110101100" => rgb <= "000110";
				when "1101110101101" => rgb <= "000110";
				when "1101110101110" => rgb <= "000110";
				when "1101110101111" => rgb <= "111111";
				when "1110000011101" => rgb <= "111111";
				when "1110000011110" => rgb <= "111111";
				when "1110000011111" => rgb <= "111111";
				when "1110000100000" => rgb <= "111111";
				when "1110000100001" => rgb <= "111111";
				when "1110000100010" => rgb <= "111111";
				when "1110000100011" => rgb <= "111111";
				when "1110000100100" => rgb <= "111111";
				when "1110000100101" => rgb <= "111111";
				when "1110000100110" => rgb <= "111111";
				when "1110000100111" => rgb <= "111111";
				when "1110000101000" => rgb <= "111111";
				when "1110000101001" => rgb <= "111111";
				when "1110000101010" => rgb <= "111111";
				when "1110000101011" => rgb <= "111111";
				when "1110000101100" => rgb <= "111111";
				when "1110000101101" => rgb <= "111111";
				when "1110000101110" => rgb <= "111111";
				when others => rgb <= "000000";
			
			end case;
		end if;
	end process;
	location <= std_logic_vector(col_idx) & std_logic_vector(row_idx);
end;